PK   �I�XX:B�]  �h    cirkitFile.json�]]�۶�+�U� ?�-n�?��L:�w�CI��V���'��� �" -�{Ѝ�8<��<�%��o������C[�U�9�7,^.>���k����rq��ӡ�Ԗ��7������*X�U�]d�"�y��(D.� J�Q�m�MPF�u-�Z���pq�����������"/�4��2�Tv�+�=��A�Fe��m,҂/���a�i�y��H�SWU�WuD<��$��$�[�-�gq
B(�!��r�"�� s�"�ED�@E��́�	�!,R2*BXddT���-�U�:��2eA��Q��I�ۊ'�J�q"!�[N�7�D2:�d�Y��2N��1�f2�J3�L�!$�P�!$�T�!$�X�!$�\�!$�`�!$�h2:����u�!Y�u�!Y &�t��¢�N����q9�$^=]�9]���]���]���]���]���]�5���תڲ�9�)���mN��G�Zl�/��q���H�a�U0���e�I�p�^��d_}��Z�PF�������+����2�@e�{ƐW��+��!�Α�.����cXva!����A�1,���\�w���!�q�\$ډ	m�`zL`p�;c�=�f;�ò��;(;�e)6v)6vPv�.,2l�2l���]X������A�1,;��<�6��S�Y��C�4�\�0pY��u��S�����6X~�O}X�:�g`~�O}�\m`�10?�1?pŁ�����gXp��U��S���WX~�O}��\}`�10?���Z\`�10?�� ?p�������B	p���U�V���\`�10?�H?p��������p�����Ss���X~�O-)�O�ߛ>r:���}ne�Kc�K#�
\�pp������
0p���`�b.rꂫ�Ҟ�M\�4^c<u���xU��-��������N�>^A:��x�����5���[NMj��Nۊ3�?1��/S�sO�r2�?1��m�7S��J����ޡP��r��-��SŜ�Pi���'>T�΂������j��k+觎�DQ����1�1�DL|��F9}B<}N:�=�'�4O�	Tn@��m�E71(�KP�>h�RN�}��Ng�ˊSw��8u�jN��c�Sw�S���>�9�����$:���I��0t*𽣢̇6�ݡ��-�H�ܔ���Yf@��C��P@�C����0u�AF ��K��9a��:�!#P�:�a�<�o�*���(�)$Hk��q��6����������;
�8�ԛ���Ի�8���$��;�8�T��ԗ��z�"������(����	��Sߺ��9�t��t��{�8�t��t����8�t��t��{�8Y���E�7��AQ�u&�7,�xQPuC!Dt_!L\���1q��D@�
F�u���
�����&���pT`\}p���0�;���x�9F_u����\q�G����W�1��:u8*0�>��nB����Q�q��Uw�D`�8�
����&��pT`\}p��@u��"��W���)���5��a���Tv���4!<,2�~J//l�GxXdl��_^�������)���5�&�a���S�yak0T��"c����`���E��O9慭��	������[�I[?e��'<,�˂���[��[?u���'<,2��>����4�%<,2�~�2/l�QxXdl��e^�̤�����˼�5M�a���S�yak0�����{ak���O]��9���.����@��E歟���V��n1@���n8@����n?@��I�nF@����nM@����aT���d�m��*&�m��fXZ!`09�o�	�0�2�3��L[EfD!4�Ŷ]+3\�0�,�m�a%���H�m��)&�h*��b��b�g��_y���i��O���ju]C]]����#�u.�fJ�+��A�����=r59������G �s�� �:�����u�0��u�fD�O�����T�*��о:��r���<#! P�F ��H��	A��z#!#Po$aꍄ �@@����7�0�FBF ��H#�8���6L�L�QH���L�L�QH���L�L�QH���L�L�QH���L�9L�QH���n�����t��t�4	a8�t��t�4	a8�t��t�4	a8�t��t܆0B���
 �#!4*���H�
���#!H���hT`\}p5	A"��BF��ꃫ�Hm2W\FB�h��Ѩ����j0�D@[y�F��W��$ڪc4*0�>��� �V�Q�q���`$�����
���#!��O��[�`��~J./lMFBpXdl=�]~�.ݚ������[��[?��&#!8,2�~J0/lMFBpXdl��a^ؚ������)ż�5	�a���S�yak2��"c�$���d$�E��OY慭�H����.���d$�E��O]慭�H����Ob~�2ݚ������[��[?u��&#!8,2�~�2/lMFBpXdl��e^ؚ�������˼�5	�a���S�yak2��"c�.sb;�H��bY�=�H��bY/=�H��bY�<�H��bY�;�H��bY[;�H ��^�&�9FB L�vG�1�`rضmh��@�0Yl�O3�H ��b�F�9FB L�v`�1�`�X`�X`�X���,�,�,�,/f����Ŭq6��`�����FBt����H���b�:	�Q^`g#!:ʋ��l$��})���| �C[4��7�r�i�cq�+7նh�š�V����ǧs��� ������ӊ�"�� gۍ��<X��q��q%d��kv���<R��N�t����5���f�y���u"���^ː�dąNQq��T�nAc"�n��l���B�q�}co��8���DN��8~��Pcr��s|���N1H���̕t�\P/��e���9m������i��Q}�yϝ"�����<���u2d �s���^ej`�!]e�%:!�|����iS���sÖǄ^A{$�C���3w dK�W�h_e��m:!�N�>��L(��pz���@Ч�jR.Oxn����?꺇W���f�</��8����V0*�C�V�Dd��ޜȂ�[�Y�!zs"2Do]NdA���ʉ,��E9���%�XH#�D�,��1��Sy �[26�I�H�� �t��x���� �t��`���� �t��H�����,��1�S�g y� y�c��T =�C�T�8s��r���1p*��r���1�o*��r���1Oo*��uE��q|��gOz7jp�&E���M��f	0�|ҿ�n��&^�F�	���Ã���`�M�^m�??,?�57�z�����9�~2��I�6���jt������� ى�g0�&^��g�����p�x�ھ|$~X~cm��j{�qx��a���׫���A��g0ʦN��Հ��:F�+`�&+l  &��"]��&�@@Lх
������!�X34YX11D�$`�&�j  &����dI��]����������0C��4Ct�fh��bb�.S�M��@@�{lt�fh��bb��S�M�@@L�T�u�n���]���,������0C�u3Ct�fh�hbb��S�MV�@@�Gјt٢�F ]��n��KF�-`�&�e �1-Sb�U�N�p��2���v��2����t��2����s�y2����r�a2���pq�I2	������9��$ j�7� � �y�mt���r���%�sl�/�e���2I8�i��џ�~L�����}��1	������9��$ j&
�N�DA��λx�����x�W�����ڼv����b��l|��aq<��X�8{�)����V:�S�_]g�cJ�+��lkl��lh<ʎ� g�#mI6g��\����`�����Ge$�"�����J��c��Ajn��1u�J	ԊtŻKm�Zv�OL�e�1S��j�T��笳_��U��K��\��W=���U�z�CttT�z�C�R���E;h����.	�	�r��x�@ިs��IݞB6P��C���R�c��&ZNn�4>�9a!�:v�z�Da�vx֧�78֧fv��y��Sfv�b��Srhgd}H�	�e�7��m�ױ>��]���l�e��������]��vj��/5I�{u�����1�q��	�P4��C�p(��áX?���P6��C�p(���hȿ����]��7��P��I��S
�_��*���ODQX��U����E��S)�u������Tj�+/[�Nsj{�@>il�y�G��2�8G�Jh���2z��bS'A,�u��A�7�$�n�F��m�u��#�_��؝�-r�}*���i��\�F��=߅�N�ݴ�]5\�� N�U�<i����K���R6��cCq�Ȭ�8wk^2�6��K�qjm�:^t�8^t]"�ֆ�QX2WĐ�5�#�H]���bD�xՂ�"2GD�;"��_6L˓`i�=	�vړ`i�?	憦'��R,�'��P,�'��P,�'����$X�O����$X�O����$X�O����I04�놈7�_N�msx�l%VB��aq��~����9��xj��'9���/�gut���ܝ�O"�մ�o� ��;~>|�y�W	����ݱ��U�kslֻ��wm��s�Vr�;��\��_���.7�s���	�ٟ7{��ö��ss��������+��OD��DȒ(�,c.�A$i2�&����3�M�`��<�e� _gu�Cm�T~v��^�!8��r�!p%w��<��u)��X�r�#��`�J����<Y�I��4~��(\��u.�ǟ�n[�u]m�r>�EA�� FB�yVY���X^�3��9��s�W� Ǜx4�T��Ғ�cdk�Ċei�lPB�j�)kC6@�'77���,�VI$�(����I�*JE>䁰5��U�B?4����*��m�gF�U�JeŐ�>�298F�X�)���6^��ZN�YOm�?A�9�o�������-��^��D��wD^���e��^�#j�V�d6^�z8�RLU	v8﷝ԟRRU��yRUe�Z�f��y�|`U���ٞ>+�[+�Y�"��j>}VM�c��,�x�>���%���Pn>W۷�e���:�������S�D��v���	������M^���],o�pP������;Dy���U��m����-���"��x^���.��o@���f�P�>w`�noo��������G�ۛ������z������Nps��i�{;��w�o�e�]��7%���������&M</i��͋CsҌډ���r���5i޽�_K��ߌ�$��K�3��5c l�&�G	4�L����&<���,9���֩�,����v�ddY�����!4G�������D����0��p�?���I7{
W?�3�f_�@��x���2��|^;G��4x9~����9zM�
L!��z�_��,C���.b�v�!GkP!���!'��B�"�݉)��Qf$F�7�LY�Ң5(�۪hZD3�eU`V�NM�hT.���UOov�}�.*�����m���,��=���2��O�V����8�sL//|����5W�^�ȑ��m���_����ܥ�3��)���2@^|�15��e��*@�Y���yU�{gkV��;��щgϻ�7ӴϜ.u]�!�8�/\�ehf�%33<�ӊEϧJ���O���9j�k&��
\�Y��|��i�$��L0�K�df;ˬ)��fW�v�/#�q���\�T���)w�bD�����o���ܟ���×����Q��N��}{�W�9�X7ms?|�^|�PK   �I�X�H<�'  �'  /   images/289c84f5-bee9-42dc-8a56-be82ea7098c8.png�'w؉PNG

   IHDR   d   3   ai�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  'IDATx��|�Օ�_չ���'稙�4���d,@`ȋ�����bl��[���5޷~k{^v��6�&�,���P	��&��z:�P�ι5-$v���Ӕ�VOW�x�ν��+�-]���}	�å�*L&��/�Y�CQu��+(**D�9�p�
�/�^g�F]�X�^7��\�-1$�:#2"��r���ũ�?���M�^�D0f���A~A�z?bI��8�1���������������|���K`���&�T/
�����D0��ǋ,�k
��"5!��"77������4q����j�"��f�ȶ;�^B��1"�!7��g
#���\�Ԧ��I�+�Q3�;r�q��������R��cn�M��@�[�!3���vy�]�H8�_��5�+��q筋q��/�Q��w����x��N`	�������133��^
Р츶a�nh�x�&�_�%Ņ���n��R�{����rMⱗ�H$X?7~t>��9���9HE��Oڑ�����Ћ�D	������044����z264y��5ؼ�<vy �����E0��x��a��������.Bw� ��,!��p��V\3�mm�~o!�Q|��e����_E@��ҲA|����և�m3 ����cA}5^~����`���wW"�L��\�N�ݠ�ݩ��أ��������$I�bg%��Dz�m܅67ؑU�9,�=���P^�b�OÜ{������>lh4���v�������,��A�[��1<�4T(Xд{=j�۰��^ܶ̌�yw"'�(t�6�Q��MZ�#��k�ȯS��t��T���>|jmrj?[��/�kf�4-���,m��So��#�H��:#	��I�9Ľ7��T�M���!�*5�Ev�]XR׃�m���V��l�21$����;s�2�+������:�K�@Sm��ҏU7K(����i~��XzO��n,�ڢ�!��+b4P�;�F$���*��fŶ��$�?Fsk�L�bHj�o:����h�v`ݚR��M���_bڗF�T��Klش7�����hlZYJ��{P����R��8?�ơm���t��K��᭽øv�'�}"�����*�zkr2Zs��8�7�������$�Y5h,����c��O��9�E���2��m�[0%t��S�8�=���?C�`��y(�t�]}X���Ic��E��q���
1DE��kV�a��q��G�ғ@na��lҨ6̯����c<Ů�$Q���X��;����F��j��˺d���>(�5x�h�0a��	��V�o�Jet����h���"(�(J
�vaӟ�c�D턂^��#ZR��Q�|�S���\;��+B:�F<�{�e�x�#Y]�|�4�#�'�R�N"�NS���<S$~G�.���PQY�g߱��SE=�5�X	���\���#/?���8�P ���T��ߩ M�fh~>�O�k�N�zS��(,,��
�z�CîD�*�_�q�;3E���D�q��4�Nbz��hP�W��4�d��'ڑ��ǳ{$Aϡ�����d1YT8�V����^"��$ɤ%	��-D�l���Q�u�e�D\V/+0�W[7�v��JJKs�^:m�B1��iD3�t0�0R�d*I�VEm�����n4%\L��)�1[�B����w�b��v<^/ȩ��~� ��j��0�%de١��$������m�98�\b�012���C�>F�!��֊90T����|���c��P>��~[Ř�f�mEg������!a�Ѹs��!|�v�:�`$NG�J�D|�����F�-��x=�ɶe���h4�i���R�:i�Gm�&BaQ�xɈDR�*�R�J̔Ĥx��	BK6�i�Äf�1��o��<���k�E���W�LAA
��Yj��G��PI�B�� U.��T�5����2�*��ܢTNՄ�.��B}:I�	Y�$ 	ڔ�T�P�L��㎯XCΟkEaI�IB��b'�:>Aİ@ ��J�見�, �2�PQ�E�7%,#W�O�\C^س$x' �	���3��H�YU���NP��C���Aj+�
"��Z���"������'�p}zz��%����R��x4I�:ю��2fn(�c�2:;;�x��##$d�}vww_���Hv��N�%$�
��X������1Ο?�ƙ�������yd��WI���b�=��J�����8>�ƈ���@5�:�?��gn0�սql��-�)d�	e�8ӕ�M��xuO��`¡�IT�¹���p����ّsIB_��w+ذo<&�"�����n���hkkGMM5IjL�l6a|l�fXbw��)ꭿn��[��Q�$SS�X�h�(��Ӄ&�{���H&j���mQ7��z���K�%��iLze��i8sq��_�Gׯ���2S�s��i�zg^{�M��o].3X��º��e�w��m�+ԁ��x��y���c�����Ļ���b2�B�԰ъ�����!a�Or٪yV�)7R�*��Nm7a��)�.@̔�+��A,u\�ޏ.w�����b��$�F���
�V�x�lLNN
)/-+~��r]�?+))���̙3�a�X�v�:ҦJɯmݲv�����L2����K�Cc�ϱ`�����<�{?U�߾�M"B��H���q��a|�{ߣ�0O>�$j���ފ/�f��f�ꖔ�����;8�Gf%\�.�@�O�MAT�)��t����,.ǯ_W���C?��*������ǫ��+
=+D�L��(;Q��_$����c/$
�`t�N�q�����C
3�&r�Ѥ�+�(͓q�3M�$in"��B+'2��fX�T�!�S����#���O#�薳-�ıfTSY;X3��O��Ts��/֎,3�k�ݾ�pG��� �FmA�ޚ7	����Ghnn�~����?�>~�B�G�]�a[|�7�����������|g�x�3�}�4����[=h�ԋ��Z{�,��7��5���P�GZ�NaIS�T�X�a�ڹ� �&2S�]��l��=tH����<����=y�1�'P�^o ���={�scppH����>1��z����\I72�ʒ���c���<g'����3	�����r!�Z�۷Oԫ���?�Go�r�ҕ9�jQ�bЈz�z�7��g��~�Y�[�/]`�`:;Hb�L�L&.Gh�����iA�X,.|EGG*+*ķ-ۆ�N#����9r���_���ĄE�2&=2V5YIs	lXex�i�/B�{_Cد~|mr�2Z�b�niFǂx�12{2z*�m_�&h�裏b�5K)|p��{� �u@���cW
{����ɕq��!	}#�4�*KPy�ʕ���H�MLkk+�4�<��9d��)Dp��f���5F��DH/�|��7#JS�D�d6�i6u�� ��,01	i���V2�m�Ol@ �6I~H �tZ'�۷4�_����W��4;F�q=}����+�C.�h��W���ݷ����sz�<����>
��8���'��&'� ��7����0I.���ygD��fs�ٰ�>nO���͖�Oߘ�
I>�/?�_�� I�L1���5��♎^N���`�N�h���,��`�;��c���E�%a
�*C�����M���eyC)-�"�8��րz��;�%p��y�gF(��OMM�s���EF���3m�4�\��K�T}���0A��!�ڋ��nF��h\B,��dԣ����b�(�C -�.J����v�CZ
��T#���l�2��.1�_W�!���p�`!�sq1��T"&a
��(��G�d/�$� �IQe1��^Mrr����h���Kv���!�h�(��K�(v1�L簖��9�9o	E�X+M�!��Ѹh�H厽F1 �L�Č*|]�h�3\Dy�a����*k��Z������ȟ����|8t��XX��Rr9+�yv�?�9ോt"M��@X��R��1_#I"�?�B�����{#I�a3bb:��2:�f��c��!���{ȅ`b�m�pd��/ፀ���1
�5�Kwm���e ��E��y+�-GR$�_e��UfH8w~��ݼk�|��.���4�.8�L�,��d��]�,B^!���	�v	"�z�J�'�q>J�*��^5M7 $��p���(|
��$[9&��u�Ւ#��/E>�6�D�Dy
Yv�Z���J�%V�b��Y�I�0)�v&)`L� ���Ե<R\�IS�0�6o��
k�8��L��@0&�2��d�/��"��-&M)���:��R	=�M:�l~��^c~G�!���O
b		�6Bm��!�xU�vZU�
���0Bg���Dff�LzZS]���#�q��?�T�a��q���W�!��)��hX��aN."����d�u���"C��-�K�!��T~6O!��rl$�DdFf�^�ǎ��mG�H��	��T6�IF{{�h''[��>gΏF�_b��߸5n&�� L�!/a�hZ�n2�V���*��bl��Z����z�Zh1iS���0�i��i�3��V�<��0�1Kuy6J
���Pt6t�H;�d��o=N�R1�2�E������I�~�̅U��뗣�Ӏ���x��b�,6tpvy�MAh@qg����NKĄ�m r1�1�pj
��$"e��Ń.�rҢT>�K�FN߳��ȯTV�!7bxx���!Z�Y/��D�\��A&�,�%|��g.�j&H(���R�T���p& �H"�Ȥx&=��wJx0l"���m�M$������,.k�10�`���db�; cb<��R�+e��R0:��#&�9�X��n���Yȝ��ՠ-��`�z뭘"l60��a{�b<#���0#d-��eM(���o*I�/�bx�S� ~��"�Fh6U�Ó��ǩY8t����J�����1"��PQ�#ߥ���bZq��j˥з� E�u��^M�t�ʅ1s?W�!ySbm���o�����8pD�{�����΋d���]3l�t�Ԣ�;�ʥ�q�zTfw��!��em*�g��ǉm�P���/�}]��H�����a�r{	Mu�l�*���Br���L����X8�x9��,-3�z̕�p��m�w�Ó*
�� f�r!c�>��M35��`H�L�/�,����,3��O@0����kVbj�=�]Q�����9}a܏�4��(�j�/�-N�_���6c�'��dBh+.�W70��#b�n�"u���n���1���Z��-~keD�^�iE~��G�$��&� ��4E����2�Tި��$��Q�d?�6f����I�K��,�KW1��i���c�P�������^��9�؉�� �֓IR)XIh�Ȧ�S�}�����B�N������d��4�n�Fqq1V�X�����MO��|B��	�ω���?�O±s!$�s��Q�PpM�G�]�Ԯ~��F�;D.�h���X����q!�P��*
�c���]���d���rƗ}�<~�u	�%B]�%�>9%����
�9����ɐI "\�K�2�'�.&���h&U��dI�V ��\a��	�����إ+�&WĹ*� ח�����@Z���		�Z��"�{�`G�J�i]�	No�+���c.C��� *st"��ۅ�-*<A�#�N*^��~��;)�PPS�mo�����3��D�,�@q�LfS>���^E���{��f�Q^����G�I����i��'vճ�����-.s�ԙ ׭)���v�X�4�����E��8Oyz�n��&Umo f�U�~1}s�}�e��r�����|��
���p�5�3���"�]L�{ǎ���5|H0M�t��L��g{�s��L�$����}�$w���e���bkl�F��]��r�'��"@u:�qg,��12��ט�V��waNyy0-��j_:p��Z0�тCy�!��9[p�|Z�R8zg�$.�:�F����g�!F��x	��% fāf^�O#?Ϲ�k�܈����!^�#�[j�z���d6� �a����TG�%|�/#���]�B�m�p�[vk!��T�ܢZ��<@�%l{���5�o\�s�SD�>�X`��gT�*��O�Zp�99��0N�p��i	��@=]籤NK�KK"h��w�q��̼+���H�g�,�s�Cx�o��{��`���I��O��
��"�9$u�0�'�-(ȵBg��e�8"�aDA����D��#?���3�$F�h�W<M1G��l�d�O���pf�/2�U��"F8J���01˾��"F��h�ef��{2)�~�z���ZD ]8�����W�y��\\�ׯ-Ś���h��׉�FFx��^�>E�����~�$���C݌����
Y���x� Ҫ��b4%�V�����*3n\mG�q'��^vtv�?;�g�
aG�*|Q�bf���y��_��� ī{�^�lY�Ӌ&2>�;?%����BE���2��؇��XVz}��H�����G�u����0k
+JO��^�$��M{';Ӣ��gڅ���P��ƀK'��r:�iS�5ق�G0%��K���1�1��5�B��fv���9�4�O�^hŖ�b*�<�hO_/:
ƀ��n�l�w8��՟&�4�=��?��bǻ�����L��}��@�9%�;���8�����x������Wط�Y$O�t�.ޑF{���'����c�Kjȇ�V�^�իW#??Oj���|������"�j>~�
�#�����C���{�	C/i��Ҳ��Cψ$�9�S���A-�sdi�u��Nk��0��4e|�u�uxі30eQ���r� �l~�z��}~4�����m����$�]���?�\I�k�A��0O���؈u�։m��6m���ƍ��؄?<�[t�]a`�[4�?�Mm��E{{Y�f���g�욅�Yջ�g�=V�g"]�Q�� ̐�����M�M��;^�m('Ʀe�J����Ua�z���O6#q�eD�:$G̈8���"�[����Y�CKJC_h}��pt	��]dg�cߴ�Vƿ>`F_4$���?���z�gp��O��&��i�|�p����?;/�u���g%�e�bzV�tb����g�XJ�|gɎFSȦg�`\���f70���iq�,@��&���S�IE�58دE�a��<֌�\6IT��XӤ�SX����������ޡX�3�S9��N
 �����_A�?C����e�#�}�s�������p�Gf��.�7�\�(�--�G��Ν�_�{?Ο�8���+ ��!,��]�51���2��&|�}�O<ׁ{�����GH��E�xis�x���8�(Ǿ�.R[3�K��up_�|�}�������܊\�	'κ�ٍ%x��v|���xys?V-�%s�FG���^�/w#�|%>�|�F�I��-��cZj��($>G�_Uu�'�.h��7$�����$p��s�����ݷ����X�S~���!L��k
hn� !��B�bf�B֋;(j<�����?,���F�x���¶�-���!���g����o�� �*�I�&N ������NP�fFQdM N��8Rnrt��#�$E��\~X�HϜ�)XD%��UM!5=M�'Nm��b+L17���.1冉ڌD�H&&>4��0��O�#/����'�Xk�re�j�̘N�bz�"����!v+���K���	$�Vd�ؑI��Lx�o^�d�fW���+�����0\��馛p��1�I���|Vd�g��;��!i\�%6�y�尀�񤄗v��΍7��I"f��Ji����E(0z�@Ll��A��X\��[�����ƅ$e�Z��qgL{v(&��m���
}��(R�����?�9{H�NiW/e��X�U5�ɦR�Z/�T/����e-�����Y[��K����.>f���f:���_��m���6�Ⳏ��J~�} �.<�"/,*��%���ZM�PRRL�������e�,��=42�`EUe	IuD�~qx���M03Y���دd#��;���Lrv=�� B��B�2`|����E�Q�Sږ�D".���8M����������"����5�k��#����(��e����(��)�̈́�y�%�N	=66*�Ysf9��*|&���˶���ӹ���b�7��6�os�1^���sZ��5��TVZ%��1e^�����	��qcaN��PaA���b�����O����9�x".���o����M���rm�Է�M�	��ʳ;[x,ٟ�ZL��:88���yb"�i��d6-��L>��&UA��eA�S�|n�	�9��eXf-+�f�)2�8U�� ���L"��Bp7�^�u����h��=����{\��1�W�&�,�	Go0!�� //�����_  ��_�c-��-�Xm%-���'�"-���B�k�5 K
{���NҚ���Ƅ�f�q����:��(�����ܪ�yP�I�F���>��<��3�u�&'�`q<����kD�������C}b�9ydBS�M@�S����Ǭ'䗄klD�e��,�TJA/IiY�(���^���`�;g7�e���O��F>�]RZ�i�W��
�1q;|0�������p�bR�C)����{p�2r�mI���/z,�@E��M�u(X�Fu7/��ۗƾd.��"�{�~	!�3I�H�$���=��Q�l%՛�ǗOc|:����W�Ҭ|�I	:���>i��˹���P�r-L긨7�J�H����2���x�x
����'ś�8��|Ԍ��+`Ӎ���Q��b@'��z��N��cid/^F�"�G��~�9�嫐k�K�8��G�*�g���W�;�zLE����2�p}Ө��n;aCY�J��q�r�����!ݗ�VA�Ɋ��6l��;�m@'�w��,�]��a����ψ|ϝ~
��eu=��xiP��n�'(��m~Gں���S��5�}_���QW���9���~O�1�o�eĵ�>���(�9�'::���6�rك��;����X2O������Rt�=�������Y������A�EO�����5(i�!�G�͟�ĺ&�l�
i`6A�'���Q��W����b�������0����[���ϑ����c'o��u7�j�6�Ͽ��{^���7c�(���Zs�$�?�w�<����t�C$�A4�}����/���	��G�&������&��Ʉ/�����$�x6q6����n�+4)����4�:�Βc�`iL���r�֞��B�ۃ�HU�T~�%��L��Թ��(��Nc{�?a@C}%�n��m��R���Yh�$s�'�����)9���f��i3�W�^
 �o��eI�<�����6F�8�&�T�pʃ������߆������!ޗe���Jh��
�k$�q2�5���>(��;dGmm>��),z�mp�	4w���o�} E���D�4�g�p��X���h�vS��R�5E�_{_C����Kho�3�9��a�<�*�Q� �"��N�U�z΅p���}��/��7����#��;VIp9@���T)�r���W���s��.���̮%I��+\��^�"�΂Δ)�����CX�����&��I��R�T��7���0C�6�63�O�ۜ8����!�d���>���(�z��^����a
12��.��`�{�=;I��z�I]9~����BJ9��e��O"�,�z�q�W�`96E4��23��_���Q.�2yA��F�sHIe��jQ�2�r�    IEND�B`�PK   �I�X�ޗԊ  �  /   images/290f8d32-1f39-4e19-80b6-a4526aa84625.png�z�PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��ipTU�Ow��`��Ȁ,��.�Ԡ�k�NY�E��b�˔U�X3�X3Z֔N���c��
��+*�,�P .D�%d%d뤷���}��N7��D�S���u�w߽��{ύs��g�-"�I
)**�X,��W����hoo�p8��M����Prss%�z�6�G"���!��c�1��X����ő4`�N���JII��L����f�����|
D����TTTHAA��m�Baij8,���{"�=�x�k�Œ r2u�q������&)..V�ɖ"FRZZZ��Ȑ!#p�`�lشY��2�X/�0JSs�,]4Y*J�ˣ�m��P$m��;ӡ�1|��ׇ��G��W����ꫯ���r���@)�I��aR���I^n�'�"Q�pR�\3k�89�2��L>�Y'�Nf��v֬Y
ʷ�~���M���1j�DbxWYY��9R�* ����⽍	?�}��pT~3{��/��b)^tB��̮��Je֏?���ژy���C0]^  'M���g�r�P(�S�ʔ	cdۮZ��q$�� �y��1�w@"y�!�' 8r�jD^^�tvv&Q��S�ʸq����������>Nsڴi
�<�~���t�@|�>ϖh+ߘ�?�{��˘������e���<�u���)Gjj%��1G��R))܄���a�]��y睧&�?���ٳg�̙3�>P-�� 2g���OdϞ=�wq]s�5I?FX�=�%+4������v�vs����-�{�>Gd��q�?ܩ�9��M�:[��8F�$�R����S=���=�����[o��+W�V��@$ �O���1c���<�w���r��* V��T�˚5k��㯯��1c�HWW�466��ŋܟ~�I.����~�A?MN��=t�` L{�\`ԨQ��ښ/>��s���;�t�_�ĢH��H ��TⱿ<��}�'�/���J�;v����* ���IO�3f��Ǐ��w�}W���z���ÕQ�}�M7�9� } <� �'�#� |�ݻw�3#F��\�(��YUU��4��8q��9 ̘h���?�\���_�W��N=d#+�Y�¦�h8$��z��$��G�kܔ&p37� ��0l�ƍ*�n�������{̽{�*3�j�I^�f�����b�x/L����7�Pf�<9Kuu��)�@`���/���zH�n�*k׮��{L߁�[Fo޼Y���K�ٱc��P�T� �ʋdA�d�4���Ѹ/��d���2��S5Sȟ���Ihe?�ɐ�;\p����Ȕ)ST��ϟ����G�������n�ɻ�� �	��袋�^�o�Q���ɓ'�o�o�������4�M��v�;Z�Y��Ga1n� �=ݎ��� �3/a���"5�T�m2ݔt�� #��ӷ퓳� �	�<��曪	0�����Y�j�j �����Ѫ?�P&L���sXh(A �AX�s�Nmk������4.\�PaӦM
Ș��>�H���
ٵk�2�=�8��G,�S�>5>%r�d8	fA���PO�+T�����/���;L˫��������K/�2��(��q	,�p|�����e˖%� 1+� 
P^L�N��I@0�j��4��t�6�dB6�wS�w��Xr�zK�e:O}����-S�{J	��N��^�ӵ���~�Ę��I�A�ޖF�7��ܹs3�� P&��s��0����\i��)�vV>��;7%{�#��f��8�;p�9�/���F�VHr��4�h�$ A��b}T����LW:�~Ƒ/��Νy,��-(í���SB/����}��
TИ�%��U�!������ 4XQ��"Î.G6��S��r��Th��I��2�16�Vh���淴\���j�C��+�"%vU;���;S��!�NH��v��6e�����Ѿ�S����&��ue�D�����+ 0�l����>���P(B8��4���w���x�Q�l���	@��N���a_�b+~+�G�.�+ �$fR�y��q��VC����2h`~�]��c�r��`�s�ȑߗ���gK��A�d�	d�n����A��Q�/1�����äj�#���V��8�+M0���Y�^��;YAS��?묳�x@p��e�r�
���t��/�ݸO��m����ӌ�k�@�D�W4�< lo?"nl��l���ΐj��l=%+��5b¢Ma.` 2ޖ��~(2���hH��=�Y{>��3V���F3�'̌�]��HT���ݕS��T-����z&Ҏ��w�:����%=�H����1�5>��>π��JgQ� �f�g��y�x�1��O'��oOD����%���L���|0�l�;0�� �E���\X[[{��� hGQ�#�5A�z�┌A����W+0���g���:�v ���b�/d.k���,)S��ws��[��r�ߚ����[O�;V�1�܈��.?��&͞�j����ĬAi��O��<۬�B'w�`�<\|��Z�a3�����M�!�źv|:8� �M��/t��)�P�DT���Y��)8���d�7�H�����[�����~^�6W�"���*9� ����=����Sc �O%DB��ě��E���$�A�Lv�p�]n��ߥ����RV�
��rb�tG��sL���,m����b�:�|�Z�)55��[U�s]׷ł�+�	L?�; �N�f��H�a��iQ6Z|��d���(=G�+b�JCm�l߱O��TB8��h���}�2U���g���jNR�Ot�ɐ��u˶Θ9�L�7u�@4����َ��u#̪f�C
��-��"O=����V��P;l�Xy���ppnKb�F"y�pm��])o9�p��w'ϧ�V?Y��m��
Ό>$���$��9�#�G���}��y睚`�%�0��F4�rS�!/��r�k���{Z�H��v����Zk�m�,��O?��^#�>�����MS�}��j(������7߬�t7�5�V`2mXrR̨��S�e��7o����LC+ ��o~�V��O?U��z)�fœk����}��^l81���>���Z`�X��m�M�<���R���;�h����k�0}��D�VB���vg��[P=˶Z�d���ZH&Zq�7h��5A�]v���܏?�X��r�h���{�-4���zg�q�q�Z�673�T@f_Z��O�5{M �瞓�M�	�����Xgo��QrM�m�&�6m��ݦQ��$��bu���cBtXl-` �l;f����K/�T���9[0g<Gf�*(L���H;��I�i��� 6��~���D����,��*(թ�rT{[__'y�i7\t�B��^;�|��x]���v�:�pPJ�a6���_}���I�=�����w���
��d��اm�E;�.]��o�]�%�/>m���֪x�{P
�3h�'"���+�$�N�AC��lդ͍��[#8���,��a��� ���K�=Y�K��u��{�>��[o�	c�(��"������o��� �@��v�Vpn�����R�e)��3�t˷-M2sB������a��(�~V �nfhS7
�����:|�����AlԱ3��2�$�9��܋���v��?Q���>߅%�sX����!���>	ˡ�v9����O�~� {:��2��bbY�,�9Zj[����M��`�}��t��Z������L�~��ѽ�3��C��@�',�}� _�j�<'�2���v���s��"���4�em=�Ś�l�n׶I&��l�g}J:��1���PM	��4vI���SO4�=��2��г_�%���gK�� a� �j^�	�މ�����Q	�������J���x�`�M{u�AՎ��p�y'�Ӹ?m�i�5y[�	RMWJ�n�q�[v7Ȣ�+d����f��PO�'��G�'MԳu�HA�!S7l��
Q\�kE&�,�Ѧ��{��4�#�>. �u�Y�G�}W';v0`�ݑ�1�.��q�r��Ps��j�x�4^��(�$0a�!���/#	ӓ��5�zs�=�A�3NT��ڤ����H1/Gj��P"�G��kAp������A���/t��    IEND�B`�PK   oI�X�<0*r�  �
 /   images/46ec3c75-1d43-4a14-938d-e2b5ecdc5822.jpg�gTSQ��B�ҋRQA��N� �BSMDDD@ �jh5�@i!JG! ґ"D���/��/�ܽ�>w���}�;3~_�J�X�\k>��?�Z9<� 8����؜|���	�H���@�����0�b�`ffbb�acg�8���w�����0A�3�.�����]��,!sQBR�@�O1s33sK�����z����`����� �5�7��X!���Os t 0����@O�'�d@���u^V������G.,��)�k%�&�+��^�L�g���\���RPTR���^�qS[GWO����]�{�v�����Xo_?� \ē��Ϟ� ē�^�NNy�������_𱴬�SEe�篍ߚ��-��{z�~�����������_][�������`��h��x8O⡣��C����;9���2riCa�/ȅ������ID�d��֫�������E�/������g@�3��a�:9a`N@�!HP��ſ���_���W���-!�H�6�\��fS�_���_�6z��:�Ф[�� 5�d{K� ����,[����/�=��x��Q����/�qxǝ�<+�0���¶f��5���N㡨���ģ����
 	���G
�
|�G��A������ߚOu+�N��QIT�5���q���!<*�|0ki��z�F��9,R�y��O�|����iK���c�R��\�ܓAMI������2o���e�u���z�́]/��P�w��/t����Kx-��3�� !��.4�QW
�;�<5��E뉦eXJ�TY�GLYB��B�.�@]T��?a�
�.�B2��� ��&��������%��� ߠ 1I)}��$�'��f�`P�ݦЋ�ʷL&�Q�
��x���3D��~#!��(��X��h��#*��fR^��WQN�+ЭQV������{���NE���K���&��\.\�y$�Bk��}�ZFm�i]
��Hh�E̜9�!j%�h��k��qeiFX��x%H-��|&n�h2�:9�dwV��?���U�#���3��{]�F���#��i��o�����6��˦~���W�6M]ָ~�.�v'��t����~�}�ה�tNP_y����J�Hl�
�i6��?Fó�5�u2<No	���G���m��Y4�����L�5���D, �R$���ʒ�sHH���8�>�o�4���u �K)��Ͻwem_����V8p�D��"k��y`u�-���f���<7c�Ժ��K�[�|=�ϑ��w��gR��n���'�EG�h�H<��Wy͆m�9oh� 	}�/� 0M�3x)m�h��Sݝ��gb��dF&En�N�`	Ա�Zf��CN'���a]
c��o�U��hd.4�>�*$E��)�d	 \� Ѭw.Y|
�����|fF3�>�Mٸ�u���_@���oXH��mX�C��>M��o��~43���Lrh�±I������{����&"B�͹/D����_��z
����\5Rx≂��Ug5Ο%ԃԬ�u1�5��n���x��,/���ե��c�g(�ꑽ���������3��2��T�t�ކ>:T[V�d���Y%����@�zJH��`\�a;��Up��*�q4���<�s�NM SS�$)rR���쟲���<���ԩûv'�e���~����=����	�=b�����(�	<�q2���5�e�Ϝ����]`�tg�q�F���UShX]:����V߁��K۲n���c@j1H~��7_Nk4�}�WA#Qf>K��0^i�?�4��$S��O9Ô�K��Q#%�?{��(t��u���yJS֬
�H��E]��s�%�du�St;$ q���%���I��,ģ��E7)@�#�
��55Z͈���@�[h�ұ�},��U�Ѣ�y�1��-��HVQ"q��5�j�I���ii��Aa��O�S�V����ߡ�(�����.B�y7sn���O�Nf������5�,�g�D;_���a~�����8�=WE��c�e��)�珱�/�K�Nl���NW�[s�� 	��2��x^b�~���)��	 ��ڠ��>i���e��-��w�"y��XJg1�Ɩh��F�3|�Ot%�HR��b���axy2֨
�i�??��%���㒦�V?��Ɂ'���w_�-1Jv~ଉ������C U'#��g���	k��*���`�c�᮸���z�	�R~�2���a����,�I�=�:��ь�\�녚ɹ_�������m@�m�0���N��
3�x�h��G���Z��ГS}��!S�y�줖�����c�U����@���3����8��ߧ"�� ��J�~�vSY�Y�5Wě����������f�lћ��,�a�u���0��_�;�s)AnN�4�8�?}L#�B�@ߺogif���Yb��x��lXG��6A2���HxS@(9䍬^TH`��p���!-�蜐����N�e�s��4��ȳ�����'&S��) Z���\������2{����aFm��_��:UX�c�#��1�߶�Iο_�W7����<�j��sXL&�;�?��b�ϾX��>��
��3�:^WT�b�	Y�q�(�����eA����JNU�������E�de
��o���1�E2����{4��@���.���q�3�	)���p��L�n|���,"�0?��lL?�HTg`}�߽:�qg��v�����;�C�R< eL���Y��E��*cf������6:�^���One�Ja&_ދ\pJ.�I���!��$�i�:Ld��FtA�^�Y.5*O�8d�K��E��ޟ�θD�&�,kI�>���1/LJ�t�_�}w�-��􁩴4ִ��;�U�q���1>���ޏ�!?_ʀ>�l�!9K�&�I�z�\��G��p�oA��U�x���D������KS��vG�h�y7����d�I�Q�7��:��`�9��P�5�0N�� �ޏ�������4c;�5�F%�����ϸB��|�m�sƭ��ԝF�R=��r��g��'� f�	1�)��S;zj�s/'5��F�v􍆬�'_�}l�O�p��Lp����JG�l�qսR�B��Y��e��SsH�f3߬4?�g�,���'�z�{�a��XTl��$�un����_���[��1n~��,�/.x���2�f�n�>SF$��@�հC�8���-_��T:3;�SIa���i^��<��^��?���߇����f�5�\���1��H�i��\ƍ<�Rp��'!��� -���*S�N}�}�l�w�V��Z[)X�d��`4v�`��赘���� ���3)����4C����h	P�/ut�
��R�)���0 ��,��; Z�گ3�K���ng�~Z��S�~O�Vu"v�����m��v���ޭ��ɲ�L���,�Q�3��`��W��B��dV��D�H�Xr�H���� o%����@ғ;J�ew��H |:���pX��\�f\���QB��δ�a*7��(ى�Q���U̯l	"�)ԗ��Gp�V���"88��'�����]��Oa��c�$N8�KV�q��@��D<���|7n��u�"L��z����ٻ���S[�,tp@}���6mZ��v���lm>�{��U�PR�.]��oN��ݺUϘ�����3�f<��o��ܼ3i�
!,!fGN�4�7y�h�<����bj���_���Mt_ �}��y���UX6���M*%����3�k�]�y��53ض �wx��4a9d^�M�®a`��4ӥL��#��&�]���(�{�fQ3c�ux@��RZO3��T�p8B���5�ܓ�3dU�;��a:q�z�G�42#Ɋ��Yə�B�r8#�m�Ww��h$<��#nL'�Z���9���q-�9ݏz<%�,�*S�D��R��N3�~
Oⵦ��vP�;��[��=��|��:�
���4W��m�VV?���v�B]���W�jj�8W�]S��o�G϶�WRN{�x���ڻ�)��ϫ�8Ϟ̫vU/�˓P;'�dhb�ς��&��b���r�'@��֫lG\G��矶���=�F�No&}A���mFS����%$��:|���u��vu���f���@�3'� N�����~q>���uaŊ��-�|�p��/7<؜^��%#w!^.�;����a+��oz���/�)���uu16G���#��@��5�}���b�-�J �!�e2O��XrNr��K�Q�H�B�e��>]켬����,p�_�g�D5�v^�� �)����ˈֈ��# ��)؏WP��?+��۰�( ���2Ô�^�2h��7\�2��|~v)�c�ex�>|ۗ`��
d����EJ�u-)~��;��,l���6qj����<�ql�1P쬬U6eՔ?{t������d�se�y"#����Ʌ�I)Mբ�g��>JЌى�&ۆ���6�u�s���>'"�w��?�:�5�������9k���/�R3`���Б)��Su贛�i�K���n��Fg�Q��l�#
�����l��!�bp�H�p�;"�3j�H��K{'+��ϵ�I�nP�^��_(�|��B�9�}����z������ٵ.0�E���#W�+TX!-u!@$'�	b	��f����h�2:�����'���*�v(�W���nT�p��9��(y��q;��Ei1(��l���>4u,� �F��.��6,���F)��^�]zDd�0�T���(w�B�C�n�VsWU����j��_�N�� (}l�'�>���42�#�-�=3����.���=B��' l��ZW��zl�|��x�)�u�O�P������LuXJ�+��r}�4O�M�ꢛ�=O�Nq�h0Kvu�)H-�����[�%�4�G`�C� �@��l��UM��)�`j-�/�2��M�1cN\�K_�D����Ү=$�0Y�ϴ�M#;��tDR�vKu�C��B��"�X[� �1��p�`��
;�Go�;�sC��9{�o3�r����y�jV�ٯ4�fV�<!a���߂��}�-�i�\��Y��*�# !��o����f*,���VN�9�{z�Dk*-�X˶�3����]�l�Rc1��np�P�}�sU�ˉN]� �IC�����zC�4�H�O�6N���'A�^����rL��5ή�Id��?֧W�����'Z:���ƫ�K?��k8�l�v�������! �?��7���i��b��XAD�3/�s[ Qx���:����C۫�ͪ��L �`�U���"�p6~�����X�@���7Nf�k��՞��XᣲiM1Ld���?
e�]��\:�ۤ�E# 0��W��囉���)��������d��c��u�T	ֿq�B@�&,�`�~��U�¿�bb�A��!3���@"�4"�y{9|Og�a�o��3�i-؁VC�th:��'ymy�vqd��Cj/n��d)3]I���쯬Ue/od���P��>x��d�1�/��z{��ea`�ʩ��t���pd�<��?2K�ș� }�3!�8oP2!���&%9�'��S��ORx�t*T�7��V?�n��.��r7�M���<��-;�@$co_�]F2��g`�Wɚ��G��Ϳ�N��[�o���L�4Ru3��D��a���TPE�:*�=q1���J��.�c�N�C���V�������xR� �OѹB������I�+��x {C��~�ňp�)R��e�X�CI��?����ջ��2�n{A�ݻ��3��)s�K�����_�U������b�āv���ʾ+9F�B�@i\�4(�@0�3���G}���t'���Yo����4�s7/�4^�Sg3߾^�We���2%Q'�(�7N�;�q/yU�!`�w�I����������a�������-��3!I�u�����S�DY^o�&�@�nс3�Lٍb,M�b�c顇��"��S�Q�s��atk��9xw}���l���Cv3gi�� �C}|u���ƈ��m�%)�h��eRAhk-)�[|M*	;j��,��a�>]|f�E�h!��9���Ο����L�q���'��H�[k±���R����?}����x\yu|yS��,������O-�!��o�#�"��'��L%s7��H고�9�P3SH�EG�$!L���a� |
ы�Fg�p����)hu���HO%�Dސm�/�5�+Y0��M|q�Z'՝���>!����Aɑ�?��W�f����B=%�^��l|�o
�$���I�� I�0vjp�;�`|��v{��j˯=΂X٨�B�u��+�1�e+|�� .�=hpc����h�X������"��s79��'y�Wʗ4tE�5r������Fr��@uet�ဇ����<��~��%9]�;Xfw���nҰ��]Q�@Z0��7�_;${b�����Mw/=��yJ}�G��m*gf"�8�Q+���Lej�<���,�lC��Ȓ�	�a�倌�,��_����	(��F���?k�����/�=b�,��N��^�L�	nQ�Kk��=z�2�b��ԛ�p���Ӫ��'|v� ��tuZ���딸ȹ5I䜧l
UE�?g-�<�?+M� G�>,����W�.����p�-9��KU�\�Y�]���o��è��z�l��{����玴?7���p���ښ��
�"��>ߠ0(z�U�f3s&��~	/`+�ڱf���
���:(���	�������v�iUm��2��$3&X �7��zδ++ �^h���U=� O��O�֞w]E�&��5BMoa��º�
i�~�.�'3�|[�p��}`�J�%$������k�c	�����~��	N�̴K[�1d�]Z�(�O6�!�*�4t�7���Y�׫d������J�7�����H�˛�t��R��y�g��k�����]��C0��%�u]�B���[��T�ɵ���D˱�g��3f���I	xq ������wG�m���Fy��_��?y�o�WMY}1.-�C���}g��n�6Y��!~�!pB���U�#��5L��8��g%��j5�-�6���n��C�Ĩ���,��w ����m���"|�P4ɿ���!Z��hT�F��:����7�QT%.�擫ND(����d'yL�/r.z��7R�]� ��lR�?���u�uV67rJ4��LJW���(�u���!�|�1-�9\�� [2��u��U�dj����k�jv�y��gqr m*���-��M%�`'�6/n���S�W���UN:{H�}1uV3=�,K�IeVm��`�����������Tw�����̬Ũ�E��	d�� ¬aW/�92������P:|H���c��/���z���?}��?L��;�p���w��a`14���>��1�Ġ�� �#K��'�t�#������n�,��nQ�N��|� ��e>4;�����=Cp��ja��j�__?���Q�� �B�r�s��:P���*H�T��7zڽ������$N�t6�2u�L�j� �x��-��U[-���
�|��5�-}��s;��{������ӌ�mA��5�y���5XUu���ٍly�Ot��/�����<@�����Ԣ�+���29�V���}��k�l=\QW�	�mH�=]�״0�rl��Ҙ��4���K�Pp��������1�c0B��t��)Lz �!P�MuT�������]��ɫ�vL�KH�m[��b��BN�c�'�پ�ϭ�z!>�{�+�ܜU�w�֒ӆ2_���qѺ:��P���p9�5&����s8R$���������u����3Ң��ʮ�mn�A�����lw^���ˡ4e��%B/�Xu��dr�6���i���1�hZ�`n����n�M� ��3b���&rf8R�D��9[ q�4h`uzCƙZ��t����]��h�`6�|UE!�:�g���ϩ��BY�'���+���EW���$�T���C�`=�6?���A������4���$c�:���/M�F����߻s��I�0PL|��;����ӌWE�h}��N��c̛xa�ʣ�%��oX���XL0g}�I`u�Wy=�au؆�
�t��S�Ǟ:y*�|!-
��x`�=�u��l�~~�ۨ����-�ﺴxj�4�7�'ŐA��`��Er;�֑���H����l��}��A>
��'��ͮ���� ������lڝ-M
��D1H����t*ym4O�mQ�͓�p��K>}�˴��.�E:�4
�uDS�2�M�J�0H���*��2�ii���eS��H�o��6[9�~0�G�l�}��vp^��&%ۇ�mr����U����A�e�M���쟔��7e|��Y���ʣ������[[/iGf�(ּu5~���IQ��R��9�X��\>��3�g�7Mr���I[T� 3s���'Tiod�Z��f����s�n�����h��F�ʨ�"2���j-�8�Δ,����X+���Â,��<� �=;��3z3\F�6�H������!؏Ԝ�9k�w�o�WG��
OWU�V9�<XSW��[�z���y)�t�E@��e�̪�(�Cg�DG�\@�KX+32rY~��,�*�=b�;�%yZ�z5���h�h����!I+Z��B��C�H[���'����L웓y�<o�U����7�tǌ��V��g�%�x_=�m�
�1�"iS��ED};MuGW� LK�z~U��|�W=�&"�-x�?C�7Q��9����<�p%�0����@�"��g�7)��!����*��j�mJ9�E���/�&��Lg����78s`7�'�.p9�,tG�F���E���E3�wg s��B�KuNd��p5��ѐ9��2 �<���z9Ƿ����0xA#�X?�x�/D(l�Ϯ���UdAtѕ,�����t� 3�xg������O{�k�Z� eBrK|����re�xw�$���������ͽ��O��?��l�wvԏ{!eSz$o��Ӕφ=c��^���\�3��D�k�!q3+ֻ���śsLC��d���T̷� �c��r$X�yX������O��ږ`�w^}�=�:}���B'��}�ÁMJ���h�z��k�u�A��r��s�������Lg�4���H<I��[�á��J/
�o����{�2dyw�ae��30�l�ty�h��q��Wwu���S�З�=��o_&B��w�\���֭������z�`N��g�_���צ}�FX�>[!KO���T�z"$����W2Z��Y�������r�ę�cutI~�2�2$��{/&�)����~���ùᛳB�:/bh���z�G]IW�
���a���4���]��%�B��xM����Dj��ߧK�V�%��>ޟ����m���܊����涫�
x�\��\�����)�����UH��k2�5���PBR�����t^��)V�n�o.�Z������t�(�%3ܬa9���f��i\
rtu�O��9�;u�š�9g'hӯ�i��Q��yH5ݗ��K���T�c`��澰�3�����Ge�h[yvq��S�'V��&%K£��'�{S����.p� ��]O�/\M�7�E����5����L�#D�:��t�mhB�u��zڡ��c�X�m��ˬs/�H(a���֡3]�ѯy��(^���!H�%0P���7Y��3U��wJ�m� .�;+U]ŀ% I�U���������oh�����ѽkx��EW�6�� ����)84�_�6��J����������x��-]09��:���A��8t����tpQ��+z��OP2f��8���1��<���&��b��Aa�@�|�������D '����1ճ&�
�U�\��&����
H�q!�:�e���'nubs2.Z� �.M���zb7E7yRh� �m4> �Uۻ�%�OL���H�Ct�u[�p`��f�O��R߳Mp�ֽ��O���b�R٤ $���1�x(1<���\�8�R�Vg%�*f}�F�������a�d��������{R�F����_���1�
Tj3B�tp�}ݣF���/ܨ}NX����ͫ̀�X�J�
*a�����O����x@�B�^�]>�~�q����?�����N��@W(�"�͎�Ѥ�i��.�1P3�¯�4(�=��SD=�$��V?����XJ�e���t�Nh���z�n,�Z'�I��h�%Ӧ2�n[�c�CU�8�tlm�e���i�����;aF�SΔ�0�j�nhP���������s��q�6�;�9�F�jh6�d }�E������;����c �O,fآ1T�?�P�j��̖�_)8�P]��{���ă}���uXk�;�H��6���?y!˿=�����1�5��u��V�G�L7�6}��|}a1U�����s��;�)�]�L0�o����^,�b?�3útr����<���Dww;��CP)e�����wu��*�JgqV��Wި�L��@݃A.�O?��)�#���u$q���x�]k=<s��l�X!�EEsv8�=���p���t^�=6�I*��5�SY�9¬D���ޤ���㬁�q�G�3-j<��Y�]��u�����%�mٴ;�L�6�K�E�[m��ǆ�ؚ�����T��w��=��U�B�P����IV�#�O�!��+YX��^��+Ю?�~aVz:�*a\��>X[�\��-����*�s��O�?K_xv���yy�Y.&%*ͽ~B`��j��%������5;I	X�b5zU��]�l�az]5��@)�튤�-wf;�[�l�{���&ک��K?�ِ��F�蒶'�ƽ@ؾ^��\0Z�CY�:���g�и۝�S���P
�h�
}#j�N<,E��,*W�*����GO�	и+j��go �|��?sVr��XD2�3����Ml��P�Ѣ^*�ɋw�93
�N���ՙu��nO��ڨ��F���������f).jl-�,�WW�!�e���#O��v;��T�$�ק_@m���R5�ņzHK#3���o�D(�l+\�y�dTj�����.�۝��搝��� ���t:���2l�cF#��҂�Su<?��DN��=mݱΩې�q}>�&��5M�G!�2���/��{_ﬡ|\�}w�@F6 !�E��!�w�]E�"N�K����W D�̥�7T�hi/ �*��1d������4�A��n�*����j4��A3jA�)L�*�]�
����r镅[��9�KG�ř���~|h��-�:����a����w-��Wa{��I�u� �(��:��a�Ƥ���'��Z��3��!�	Q�Y�Q�]���L��Ͽ��o�c�*������H�_��Esi�馐�!;�3��ɥi��_�ߍ'�9|.�s�8�9������dK�@pW����<�����}��'��p�6����Ew�{�����Q��������Z\+9q���*[o0��>� �c��@��<��z�N�YtT��~��gtb� 0e�x�E�J&���|���0L߅���|�V���uo�3`�� ��0�˷Z�:�*��g1�U��U�]C ^����p=і�$;B�����<K2���P
��g��#�9�6zd\�d�p���r���h���E+ꏑƫ�[����3��c����9����y\8l��HgVI�A���3E��a�1p{8��U���gu`�:�5�ō#���կ��^\]��(-��0g[W�t�ܞ@���nqIw�^�(�SؐY��2殛�����o<bv��_]S�8#ڊR��b�݇�Dβn�c IY��(������nR�K-p}�,��������e������X�t�#X6�Q��P;g6���=5������T�R���j���½�M�|!7��*vH���Hc�eOt�.�dU��W7�&�]$�p�gGw�-��L:e��8�0���W7jl/�*A(h����b�KQ<1�x�Pz�s�����i��{<̼��5q�σ��9�Ų[�s���U�}S��gwt��,�*��D��M5�"�E_�gf������
�DT�D�O/ГW�O��ڙы�\��:�>����&�R(;��ۜ�h�z&��W��'�'%-F�A$g��j3���Q"ifl�����L���8����D����R��SGu\��}���,���B�����4�G<D��`o�'S��ϫ��=n���R L�͙�s��V�eo�j��;d���O��
8�1��Փ�_�#mW�E�zA@��$J���3�6�T�U��b��C�u"����ؐ��Ｐ�� +#�
�'uc���8nJ���8�����PG��z�6*W\]�Z�8�g�ש�ǟ��'�^�(��t!h��9<�R{��;�#�FkKwi0:-�쩵=m'�����8B��x@˖!�g�r��n���=ګ�3%�u=}�[n�U����sl���L�����H�w�:ɽS&2��'�a��g���/��������{�L���-��B��H���)����ɶ�v��[����cVG���@�C�'K��9f*}�D(@ݹ}�I���r��Hň���b>�ŀӦ2���u�s�
�j �ay�"�[�j{c|ZpG�Sɬ"���ibE�6ρvd�b[�)|4�*�KG�Z0W<:xƳ�s&҈G<ّ��)��\t���G�LJ~[�=�lT�� �';O��*esY	�ʉW�d�T�g�Cl(�l��N�d
wDZ�O `ח�m�UGg%ND�e�k/ Oaw��-Z͸�E�|z#:��C�[�ֱ
��ő�z�<i�j�r:�ْ����8^�/��@���ci&3�Z���hS]�܁)��ڵP}�ֆ��V��NE�/�����&#b�F5r��½�!�e]^:�৛>̞ATVՒs����[}�@����Ƶ;`���=q�lj��,�t���w�eȕ�2���>u1)K�i���a�Lt��G���,����?��b=tN�eZ\N�=�sȽ�u��v�Pq�8�}��$�Z�䫲~��:(L�a��XƣvvÇ=��o��˙�/ʞ�l�N���(���	[�u�xݴ~����+�B?����)���o�.?�Щxu�^�˴��<xل�/������,�E����K"�`�Q5SG��5�
JѯV��녫�`ـO��eP���/��Ib���'c�~Z`�CF�Q��y"`G��}��g�D��z����j軔�{��0�y���� |3"��z�3��U-����4���\_1�O���]���)��ˆ������s�V���?�0�M��±'��]��w~$����`�^�*�"^��p�Ǔ��̂h^AR-#)��,�M��e��� ��Tq���\U+�6MX��=��q䟕}x-���(<�T��l>B/�aɝ3��GvJ�yC���?�G����-5��&�mʟ0��	7��l
=��H�������T�_�]>E�A��WY�^�LDCZ��+����� V��{��p�-~���Ħ{�*�8�g$�b�h��-�����^�i��/�k��/(	fk�_�~����a���3��a+e;�����l�Æj�cL`�8OE���EDq�1� �f7�*���+ĪBWwzby"[�=)���K�}��4�Ym�Ԅ��fDg�v$*���d6�J�˗ѫo������ ���:]w��K�A ��he���F�ӯ+|�]]��{l��H���P� k�h�&�]���(ku��0~(?�J�#Z�<���k��!�#��O��'S}+��]ED�����P#����)� @�,0��$��v��]6@��y&dfK����1�$�v��Nu0�{\C����_��_Rw�aZNr��b�[�1�ztb�óZ���� c��b3	����O%�'���֊a���᠂2DhN�e��@K���^����v'B6���� �.��o�y�zR��)��
e�U�e΍�7}W�hVW�af��I1��ZM�k��X���F8T�8�P;�����7���"����.�����Qؒ._HY��^PƼ�����=B[��)�x#}7|�#t�qá��w�����	1f���̮'Ι���p
�}��hϮ��	�9к9�SzI���^]���������hf[v��׺u^h�gC�S�����a���?M>&_��E\�f'-�/Rn�'����fY�|
���zX���:�-,狊�cBuu8���Ɔs$��H!*WLJ�a3f��Tͧj�M�G��鷠]�����z��@�Bj�0�\�ui��R�M��u��_rIV��v��c��o���;}���/yF�
,�[�����=c���`.a3��P:68�Y�����s�?���L��Y��A��ujn��1[��~�����Ha�����7A||/w���ŉ�����?mm��P��RL٢!A�P��`��C�E���O�|��n��Zd)9��f�։u?5�����le#d�{o��v���z�(|�:�P*����cچ��*q�4���z�g��\�48�d�}��=�#���4ݽ��f�<Y{���[ҠXC�D#=�8���u4�,p�~9h��R��s����V���9���j=�X����ۼ=����o�ib��ary�3H�̀	6�U���G�����BI�P?І'Ԝ��[�åө.jaeow�']^>-�����C[� 'T��ϓ<n��9=!���D��K`����S�	���h���v;�{+��4e,+�}	�"���2p�9��`�^�İ�Hat��4��gC�a��W�z��b�ɢ�Z/�K�p�M���n�����B�T�¶�c��:�:Z��fL4+���׶o�mw*^[|?��]����T���Tq�����L����|T.D���[Ƴ�ik(�e�9]>^��#��"��� �ԒI��N5����t��A�oiVeva\
շ:�%C�!���ϔ|�PU��|
�ޜ��T- $�F@/�7*i63�a�x�)AN�Ea)�Xae	\O3���y�`�xK��d��8�� '�~ͩ��ؤ�����uH,��58��z`=xp�5��N�x-?U�D��H?r�~M�\�9�!W0�R-��(Ͽ`��J�Gc���B�� 0ל���uro��G7`�o�>�p]|oH^$�$�r��ؐ��1�O1��<$=0g�AE.D �XÖ9�g|��L��Q	�5]���Z�0�N.�[t�]	��u(ѯZ�﫡5�k��r�z߬�i�89��@`�nfl�ӊ�������v{L.����/܎`S�0z������mG��3��|�:q���Se��ҝ�x����ߤ�}g�pw���+����rZ#?B2N���E??�{�(?����X����kW_��+�o����#�|����&���Y���6/r��ܜ���w�H��H�p��l6T3Ղ\bQ����v^����0����L�������Mԑ?+��:8eÒC����Y(�)O�Q����ۿc�L�e���+b�F9Dg�#�ȧf�ﶣ�� ��Ɣ��hV�SB[z�p��V�ӽ�[~O���P�#L�6���R0�G��a��	���8�\�挴�6�)��<
��N[�reIO���pG�	�W?M���z��\B�p}f�9e�)��5�S��?��+jDū�}��kl�M\������Z��g���,��9�w�P%��q��é�#���������̓��0-E��uʷk�.6���5r?,�p9�������r��� m������u_7'��-E_�Pu��j��������y���c@u�;X]aL���%�p���#�ɇ�;EK�#J+�Rj���PDN���w>�>�F���sHk��@|,���x%W�l�9�������=���7��w.�8\h[ `�&A����y4�uф���S8B�`$nG}���I��Ù���ߐ��.tۿ;�/2q6�ye֘D�"�f�lT:�>��~��r��叛Gm<p�~1�~��`쁿�;�f��o�q&���[b�At�l�g��+�w���^8>L�^q�]�"�*R�N���E���w�a�B8ry���.�.�٣�J�c:ӗ��qx"�t텫Nr熦�������]tq�>Y�|2_�޻��K����׼�aԞ|+�K�/_?~���ԉwN������<�m|R�e-�[(����܄����@����3����� �)AA�H�	PzW���iJ��EP�W��(]�Hｉt��{@J���9sg�3�����b�d���g��}�S����P7$н.�%� 	�T�]� + [#����:�s9=(<���,z8��$�������Dݶ˲�d1aR�� t��A_����ј�F�u3���j��V�U�{� P�<�����k��)wc�^Ġ��괃/�Ot��C��5�?T�쥞E�0�@���ͤ���Ƹ��l����ΣC�^�=z���%���(ᵂfB9�[ă�/oX#ډ�d�u������(�P�����J�2��'q�O�O�����`�����I-m����΀dCMp��}!�1�9�lP��
�DQ�iyN�/=���C��
o��z��`�1/���a\ƳH	�W�qJ�@�J���7G�7���Uk��������T[��-J|YK;��Ǿ��z�ĉ�c	lR-�R$��Id,6��ԅ��W<!�%>b��"��qS��C�;I�#��\)]#�-�BT�����DDR��vPm�q�dn&��A���:�O���5�y`�6�k����y��ߥ��sA\`��x�W+�VX�\�6C������{7�����N5<��ƞD/�]\��������i�z���d�]��XOa�9ꨜQH~ �Z��_ܼxI��v���6�W��w}g�Ub�zi�\$�ؙ�Tx]EK�+�c���˾��z��i_N������<����ڦ���)�-�47KO�}6�gH6��15�m��"�k7˝0�=�{��YމfFdC5�㓢����-x����)���{��+*r�M3>���0��4��K�[a�.ｊ�qO��k
l_v�����F^���8��e�Kr^ٮC�D��1�Lr�c���� j��\���2��%�8������I�3����ݩ�Mi�N���B���C*��"�a)~ʳ�5\'��h�[:�i�e(�*����"=�}���&��������Z��"+}3�ܻL`���FN�_�
R<�Hl�Ǽjڕ[��,}T�,_u�L;8=~�8��t��0b�S�K�~	B��V�X��J'�U"g?i'����,[i\�����8UǛB�ӫh��M����c8�4W����G���E�v��;���:��.h?n�P�{t	�ד�ч��_�,(��.���}��O�n0=-{���
�Vړ��]�z�ڧiJ��iOl�������o��gp0�)�^��4:)��4^G�Ύ`"w��%�Y=��!N:��-�)#=�d�6�'��ARzG�@�k���i5���`T����V�Zߪ��T��h�FN���մ�w��gqq�U���7��T��d�	U��n�>e�@���/h��oSߗU5"��K\�P=��+�C��'�����A�,��дp_$���u�:vUG��􀚵��Jƕ�����.lA��=�g�蹩Oes�.���BAB�A[�&�)��lE��9���)#3�^4��8��1:T�VI���Ӂ��V�����h���$����ܧ�p��^��p�~��~�nsT��CoX�'۽a�g&���_C��=��n 6W&˲6k��off������Z���E��S\�-�v�7MV���6鼎EM^��e��<�'�@��΅��6'��2�oo��n �����?q��7+rT_sg�$��t�9�Mֱ�~�&_�*
�]�u�zK�o|5�j����V�m��Ղ�*	�ߵ?*��jO/�]8.�8[���b������AH�;"?-"�t����#�6ȭyI���wS�ruSk���kއh% iVQ�9�o"`�nsn�ċ�:��"����'H�荴WgI,@��1�:�O�����	\1���6[S�A	³�B���w�e�h �q�ي����c��(('�пW8��s���!���{�-ch��ԓh�i��f�6��h�a���@,Fz��`͕�6��2$��f���M�n���E�,G[���D��SږI�a�����D��GK��r�:덴It�)��D�ԯ�eS^�g����X�~�;�|	C8�ɇnTA>���C�6/6�A�_���4��"��Y�Eu�����$��+]����ۣҬ.�N�";��jg{���O�W�ls_��(~|-�'i=�4xs��v������;X�jt�O�+��<�~�4�9���[:Pq�&������}�M$��6�g�|Q��z�"�t���q@��B�8��xn,u����� ��������},T��6�K���c����S����L�7������@�����w� Ə�JB���g��/�PT.��0�L� ���3F��_�`��W+M5Ac�S��F�z.H��=/u�S��\vY�-��93B��"[��t\]��*�Q��z	�7�D/�u�?&���s-�/���)	�[�0�Yʛ�V��D�\���]q��ß�H�1p�u��)����i��U���4�x��Hφ�y�F��*(xj���ὂ?��\��:Im�u%a�{y��)u �=G��3;۸/�#�y��D���z�M�v��4��p=�;�It(A�&Tǡ�^��DO�k~u@(v�N*;֔{���b�6s�%o�����1S�(� }�y�=^(
��K��$�3���W�^�]��㶌���c~"#!���a���j����gl0��')Ğ�ٻ�)L2Ǵ������L��gP�����_4%�İn����9���;Nn>�7���\h����|������^��!!-�w�[���ŧ�|~����._Wb�R2!��e$[��D���B|#��N���z�l��ww/���Z`�����6�C
�/��Q�A�G�Q����GR�c�*|z��Ip�f�oG�TGYy@��}!/KD|׼��t��l��.K�b�{/�F�Mn~.쓫�cƣs[P	�3m���)�D����v ]ܪތ��9�Ƞ�@��ﳫk������>�����	�E�~^���E�=f��ע�4�;�sl���1E���,B�}SN���-�D��dq�>\�T�.�d?|ͷQ��1�eQτ5�գdN�}��7O��z�>��(�\�+Fϯ��?Xn!���^e|��Q���˛��G}����F��`�2MAG�C�A瑀��Jp�D��{]���uӺ�@������Ϫ�V���oY���C>�HE�|��G�<�>Th���F�B���@��_\͡��S	���Q�6X��ϧ�>�>yT喧A����%@DTB�CD̳�M:�O,oud�͔֤]ץŢ2�3	ݚ��请�/
�`*�AM��oHTl�"F�^x��t����|�ʢ	�S�E������&��{�jR��RF�����w�u7m�{��Kϖ!?P�&hz��� �ɻ������/�2���$[��������O������Kp�����Tb�g�ޘݯ����,c)ŋm�V������VtO�%�8����(�u��x5m����ϋr�h�zhє�����ί�����DYǫ�/{J�4g>_������͇��h�03�5���S�k�/.�W�|��Fsk= �x�@g�s��^H��L��<�|��>Ǒ~�.1�}�O$B/s�Z���`3�ڏ��e���O�'c�EYNbk%�<��n����8�5�fl�'�ݓŝ���(�W�� (����w�1HD�U3VD�:k��Kz�X �Iʣ�Q1_o��?�0��E�l,�l�mC|��o�����]���v�O7
-�`ۘ�����棅]�d��l���__��~l&�� Q����t���2���Qm�?�x+j{.7�ZD-z�otZe �qXq
2f8Zm�	K<3
����=V�8T^63*��B����S�]4^d*UT4�j+a� ���C���5�+�g�wO���>��|���p�$J����H����KSw�i%Y�v �� j� �#�Y�]h�JKX;���^�YL��5�inĭ���7Ż�B
��eލohzg\�x�f��*�DN��r��I{ݝ?~W���{���ZmQx���q�{I�i�N4�����?[p$��d�M�%�ApjY�ߩ.���q�,<k�踡�6�C��Vbp��H�񼕔��\�Ҩpm="���**:ڹ	����$={���);E���fתj;+y�A'�
��d�ɗ�PYW�\D��O���o��+Rm~�f�p������Տ~���}a��K�/u!/��K0 ����D�"���Y�<CJ��0��^��`�ojM������8�Ln,����f,���t��V �G`B:J����Y�d����/�
�n��|i:6	��"ʣ_�y	Љ��s����!SDɾX�6���w�^��������Ǣ ���	�}��B[�vv��J��qs��[V�F�GA%��D���W�w������y��Q{h��==�����M���]}��(Ն�<t�1�O�2�}/ q;�Agv���ZZLY���N�r��U��d��
��~�P����Sci�^�1�];Tu}]���PEz僽�X�4�̋'܇�M0���i�ء���]�5�_�6�����nmP�d�.��^�
x�}Q{_�-��S��<G,W�G_�Ȫ����X��c�_���z��E�C�3����%���%[?kE�FfI�˯?n�w0��d�� �]�R�=�i�Y� �S�e�7�:����n����m����h�	V��U��V.>��.�7��T��;A��-�2��1қȷ���T����b��~��&$�W�Wy	O���Z e�X(�S�׃���3/��k��qp|rab��2�g��ȑ�:�w�/�YW:���`a���^}�ֈ��Kve'Z��3��vY�z�>-Uk����RZʩ��[��g�Sf;�L��+���ް���gI���9\�����(�l�`��k��1�,Wo��T"�������Iq j��h)Ɓ
	Np���D ]K�!�J�jC5�a�v���7�� ĸ(����Ӫ��.67SE��_!�����Fn&�G(�VVa����˺g{� �m�������IEو�k�ʁ�3�B��;��V���&G�����ս�uS��jE�������Y1ݒ�엋Įr�hR��I`����)�:�TG�m�2�f`����4h���EB߳�%~��2l�e�*𙹠��*�ӯ��!d���t��<KR�����'^�Wa�`�-�V㵽�τ��ԏ\]V^ɨ�˃g�_S�s�s���M�p��Oi�[�	_-a���')�����J�w����/��j8Wc��p�o�B�碥�a$�N޾��M�7��X�%i~N�GW���7��?�j���7�rT��OC����xeۋ�H\ƛ_��~4�"��#*��9gN��Y~��FD/���u�[ZDE���
k��D��'.	E�,��(]��@����=��*��$b;�P�a̙�yo{n�t��|!NE���W.n\��LXW<5�)�p0hnΉ�uнiR45T� |��n�Kp��,,pD��K]�%��u�m��>b��۞&�.c��V��Ni������x�r2H��j���A�$�v��Px&,0�R����d�D�o��o �B�k^W��.b�.Ӈy�.QC�T��L��MY/�J�S��u	>����s������_�D<?��r7�����L���L�dW�wE/�'en�q��=�щsK �/��ԁ\C@��3���X������hּvf�@,� g�U��K�� �^�Ԛ����v��5��ab�L�W1�n�����x�.��צ��.��ʳ��=�}DT�7%ǝu�ju����þ)�����<<��aK -��8ז{/vV7�kx]۔����]�od9�{�cZJĢ(A޼�d�,f�O�gIv��ۂ
%�i�+�P{d�'�,�z��4��o~U4k�-��)`{K��5b��.�f�����I���J���Q��l;�4�@[T�܂���0|�GyN��I*�������O-В�n��jOW>{���dne�č�W����y�5X*m��'��?������l8|?�(Q��f-���Z�@ ��x<[��C�לB_.2�<�<��D��%C�C��rwdǐ�ƶ%�/��p���ʒ������e<�hr)	Dƈ����{�*�\�K�:ޓ��wC�upʓYL�=�Np�� .��'8�f%�k�K�9��u���N�����:�7lV���/.��^��Z%��N��9v&oZ��䛚�Qd�A� ��wE�Ľ|_yNq������o�SI��z��%F�bj�M�,�WJ��^H���zd�hS��:"�k�gҔ/�q�]�aY@�q�� K^H�rػ����㰗k�o�a�w��[	���6���nߪ�˃	��C,�xBW=)��˼;�(���Ԃ���Ī7�{3V�lb�8U�AJ�}a����Ot��C�4;IJd���B�_ ��&�~�lR�/ʇAhB0%pv��K{�kǂ<�g7�)ҋ����u'���嬛*?��Ĕ�]���W�2���0N?+`����d���+�@c�b���G�8�<Z	�C$}yí���UT����'�QLk�*d6u��O��bE�G�9U�ĉ�A������Z��Ũ��M�\�l�[�|1�'�"����=��cs��?	m9��u�{8�5�Vg�}[p��B8p�G^vz�����/��Ƽ��Ϸ7���Q�::{:0�$�� 4P�h����Z��X���Z5k},)�� �[�������-��Sb���p�w�
�J���Y�p��m��1�bA��"i3��͞���<�9ϰ���46�;�M��_�!kw+���Re.�"��C�5o!�zYKz±Pd����P$r���U౺kǸt:�pKg���S�#T�q���Ze���z&%�4�?ٕ�4T�	���nJn�=��K����ˏi�$�&�k��-Q�P��~(��/���މT���75�SK��f��o�$�����R�>%1'㕈�h���B�����aBv�░�]�f�F���C�m�[=�j5����󁚝���)��-�`/��˺���y��|x>U{o��-ϵ�U�2l6�4�u������V�W�螵���0k9�VX��,"lq=#Qp'� N�=@*�����Ԏ3I�b�#�,~4~z���KP>�sSq�z^،T�N;썫8�[���Fx�]�,cc@�c�5[�2�Sx]N�v�-[>�5���-���ܟ�q�2��
|+�"+@�6n���Υ�{Uq+�"���p@�x�h��� E]�䴝U���U�n�KJ3��'���p�.3�h�n�ՠP�|%L� ��4x��:�0�t_[�Z_|S>ҍ�M m�n�ݾ?���F�Prl��K��7�li�S�7Q�����_� /��ṽ锦/U����F����{L]%oY>�<�,��S̈́�)ޙ���Й|���;���}�8�ш"��:�du]iE��g���p�W���s�?�,�
B�cYh#���X�|��N��v�P�u�� 8)N�!�S�w�fl�:s�gg?� v���j.�/	;6�߬|�00�2D�C�z?Z4��E_��>�?D!��2��9��V|ߒ���~ӼP?�;�i ����M5�;��O^dڟ4��v��;�;�<(d�Ю���*�*���� �����=m���_ק���U$�Y(�Rp�����i;q>�
9hv˨�XӖ�(>>9����i���O�%xX@�c�Q*�*7��	�J�c>Oj�$�(��le�~�Q+v���������檲_��n���I��yt�q�r/��bޑ��|������u�/?�H���*D�VM*G2ٻl�V���%P�d��q�)m��g�[;ܽ�W��{d
-�V�������c���&;<�bKɆ�>^�Ѯڷ=�5Q�C�w��L���!C��}>;�y�'��|�Eox��b)�G�7U��9�����Y北�5Ƌ������T��
V���X���4
n49�Ld����!��S�J �ޟ��*�h�|�$L%|=�.��n/���m�/E��S����;f}��ʈ!<-&��(���{M�G�0=�a�ƱB��fM�1��V4����"����;̒S�s�f.3��i-B0|y{�Ѭ3?k�4��L˓��!o�]��_�t���#����Ю�<�N�s�@�hU[c�"'����k����Ot5P�ֳ/t�m_���S�ĩ@�!��:о>�[0��}����s��:MW5K���>4,�]�nD۲RVL�8*�͕�眯�Q����Ebԯ�^Zg���,��O���6]��m��;L��M��h�1�G+"Y��%z����F��F�}��geAӄ�<� ъ��S�����u��͛��?A�H��9x���D5�_����:�Y�% X.%���Ě]x��ыG�t�����-R�C/��ƚ>�:^S$�)�a=���O�
�]�̠gנ�q	T"g��#ă�Fu�r�g��A�=v�<���������_v�f�+db$�ukDv./���N���A��g��Sp�9�z��m��(h#~RR��_���$��XW[ą����a���r4�Y,�o�A�NK��!h�q�:���x���鳍$o��;�泉�pD�JR�]=���>:�VQ����ob�Y��Ph!^��Ҏ��V���7�xn:�К,�/���N[��i_�
�Tʌ�\�1�OL�Ѷ.��cSN�iT�����p�3~i6]e�^qh'�ߎ����	`��XHSkr�Q�� Yy7GY��.G��K�	�냮S�4{C�Y{	/�/],�"��Q�u_��ւ�=���b��Y�ڢ��v��3jR:�.\1%e�� �!P����.ZO�-�KB��:��PH.��D�֎8Y�7�kscj�����@ho��|�*�`b��!"����Rv45�юl�`�P���b�ZcU[�I��I ��_2�6y3
�_
�`�����8�����(ۖ������a��"�=�..����?eC�sբ�B5/��r��!H�?�˕3S�ȽG���;J���{��VC-��L# {9_�ٍ�)=���&y�}F���ߎ�ݕ&$&*D�<}.5_����t�u��My����:k�3�n�f����/		C�|7���q4$
mـq�fS5zz�h��)�'�Sm���e�u_�/O�����z3>%�J��˲38��tU��Va*1�rL?<�3�%�~���g ���-��s	��dS%�x���&15"x�.�1�Rݡ�W�����a��(���<Ǭ�W�߫��yUG�/�f���Q����g6���~��|s�CjG�B�b2�۰r�$��a���<䟠TʘM
�kzw,���yד��L,�j}L��YI�F�Yp��b��l���p��m����r���U�=�,<(�;��C��� ���M㙙��2�3x՝�uHmL3�k��j�1��p=�@q��i{��C5pH�g�T}��.�iA��u7�������q=��jK�`�Nb9����#�۟�������=`N�
Z��dν �w�{�%��%�2@���_($�V��>w:�8君}w����T�O1m;Mp�����翡|a�vλ$�:��zH��U�*��� tT�Ƽۿ���^*T��T��v��B3sT���7���5�}�%�<��Z���T���NF�RE�<[F�y���~2��R>��__X�l*s9�Cg�� �bda����;�K��!�$~���	��@�s�7��������K�o-����������_��o�륜r�����P����^��l�PWA��|H�=��]V�y�i-�r�E8� ��W���Kb)�a��G9I�X��Ѝ��Sp�-���T��?yǞ(H�ˌE5�������a��5!���}�j��x%�����?�E�D1�(��<���gÔ��~Mh��%P�m�i����	�о���U������"7Pܔn�"ܛyv���)�E9v���OLN�o��$	a�8-rN̜��x�_���v�b�F������bǅ���v�Lrr�H�E�k�2U#�%S�����&�-�><Ф�N��GֺX�P'�A:�(�}�華�m`���|�M�pV7���{��C���*z��ײRU�|ߡ�r�0}�>�.�!!�Љ�:o2=	YM_.!�i�o��k��gvm�ע�~o0�jn��TB$�X�z��lz%������Y�@��;�CY�r�m����9j�5%���ɞ�_ߌa!,�},7q�e*
_9S���(�Ĝ.����"�ѱٿ��#���:C,�X+�|�֣rC��|���=4U�Z�h߽ ��D#�i���u�Oz�(�\tt���2��=.�V��{��j�c[ڛ����jU_�x�%Yl�K��J�SQ	5��,Q.��D>]�L��5�d?�s� �z�p�|S�!�%s�f��3�/ࡩp����i�߾)���G�@����F��JsW�M����d���L �tOw`�Ť?;���BTda��5tp�Ġ�c�����B��Ņ�t \C���$�	�����1�ٝ��U���Hr�rG�Im8j�լ�i,ES��*��|΂�b �p�ޑl9�-H�CYj��9��,��z~�(�<c[�_�?�m��<�k�y|�~���������&���\g��zN,բ�]��4���V�>�Y#Z\��*ח)Ҡ��3��XM��YK;@2�f����Q۩����^{��sс��x�-�b���8G�R� ���b�@I�������y�0���^��<:5�[�D�וEC��TD!�~�����Õ�-om\�O���-�*7���2��U
F��l*�ۦ�W\h�S�Q��"��͸�D����R?J����I�p�"*'���z�R���ܬ�K��|����w�3$O�м���R��3|���_oS��~0.��҇���l�%�t
�ض�9��z3R1��F�}	��|jO���X̝���
���	C��QȬ�i�hߑg��L�l8[��H��0�L끶���jn%�)�M�K0�K��O�Mc���_:�4H���݋뚢5=p|&M���N����׵�u������;_��<ЦXq|��`�!��_r��*�S�؃Ne�/9vf�J-�� N<��_�`
{��X�rU�7����T���_K��cg8b�ʮ8���6����>�����*�-yq7̀`��Ծ��\%7��Ok��>�W�C���Ԧ<!�4�1�|P~�?�7U�pK�1�4ڙ�M�H
�nF�^5ɟ������^���8�B�˿�ddާ(�e_:x����BS��=lj�/���RL"�:[1����4_Q��9�
y?�fe�P�I�~��׸;O;�~|���?͠�_�����_S��0ѿqs��<:.��#�l�+��k�]俧1':]F�B;}?�iO��M��K�5���p�����)���ə���"�N�zf���Ur?�wF�E�{Ӎ$u�!�\��]6U�骻̲o�,ʥ,����7b��|�f�Լ�L�T:g9>�F�'*���v�qj��yţ��~�;�tQs�e��ɖs���b��
O3R���V���qkiD��b��W,� �����X[hV����
���З�Z78�F^�u[x��o���'�[l>���Ř�\T^��b8��tW��K�Z��xؐ/�K�~����vm�a7��k�ŻAR��[�a
5��V�e�%pM=�zhu����!�r�?ȟ�g�#C�)���nߌ�vu}�N�7Va�8���9i��Y̠�&-*3�p���b��H�C&�u�.���� ��S��ka��}RR�����C�ܨ��i�KF"�\#�c� x��y�N+�w�p�gWfq�]�彘���d���+IC������i���z��L��S� j7�򷠨z���Z���R�C>�+o(y���Y�豕�R}�<�2U$��k�@X���)��f���� ���#b^m��:��.��1��v&P :���%�G�̢��>��}3����%�Z,���8�Y��6M�>@�~��y�-W��t*����ǉA?Iګ߭�h�" ���Ʒ`֒��� L�����`�%���!�~w�zO��M:�(9��!�+{ "��]��[�b�4V��c�v�%�2�jHt�OxiV�	K<�b�nG_�gY��nt�-��+���.O��mhsec�Be�d��e��}�Z�����g@	��I������i�s�F��%�*��I��U߃�CFX�GBQ���B�?_!�p��Lڝ�vL�aO���-�_�x.�G?�3!�oa��\I�IUa�Չ�w�����n�H���"�^�-g\7	�@����֏��Zv-�}x���K�����V�\��]���ڦ2�8��Yy@��K�"�-ߣ���> 2�q'Er�{]�7���,
�h�/|�� �H��j��vgS�xg�3��b�����Za���6fvLg�Uj
�����t!�E���l�/c�f�G��voY���N�A`�S��M�7+�y�K YN����)�����r�;�L=�w��v�[��]cY�$��X���Y�q~�h���1�C7�v��a򳼩��k�����^�rYP�t�p�����)�{���cs��b%ju0ꁥ�/�Q���ǒ怈EmTV!�oY�#����|1�~���.cJ��{Ȉ��o��� �b���J��\Zei_~��{_vd�[�i�8,Y�����"��W]��аǌ��n��q?影�ں5M���m;|�>�A"����7����&{��>�Ub߆ � w�7���A)������	k�$�U�=R�=�br�x}�����N���VTb����CUskc�5��{���|y?�M�+�m��S��\��q�i���.底�׵�V�M�n��e��pA�8�<���������?�<��Qf�{j���X��N��i�:}�Ï`��������;�?X�7�a�������9nZ�\Qy���BY�P�ˈg��쮤+k|Cp�9����F�r"[{���S|	%�m�ה��^�%������8�Z��eޒi����>����<盇��Z3]����<��;mk��f�����TD��Ԃ4��[��)~�^ZiY�9�[u	��H��'{[�u�T6-wQE^y�u5�c_�VY��FR2�Y\A@yڨĵo�5̃?p��Q!U��+�"�!�~�=5���5ҝ:1~�ȭ8JQ�_Sb���q+���IN#ӣ�ERg$q͒�i�	Ǐ���#���x��B��ϋ%�&�\�?���RO�5QO\�*TDD��r�];��c�}��J���c���+�KC$�>�H�m�����k���S9��h��qܣ4�S�B��^h�P�}o�K�H���۩e�)B����ql��U,u�z���/_�'�Jk%�䙤)��U�=a��5J:���E��Ò�\�[$M��<��_mg�B�Ƽ3u�V�vT��G�f�Di�I/X�pĹ�`�9 �GBq.��Re�o:��l���ƣ۝��᤹�*=�E $ͭ�!�%��>���r��1ѦvF�v�in���8�l�n����B�K�� �@䫘G���'C>K�Bk�� �\��X���H&#���抅s%�4o�B$G@R��r 7o!fq'��Pn��#-�ζ�i_�y���mNa�<PC 3���N�Q��+��E%���r�����(��d4@�>�  jn,g
�yt�p@����wr��'AZ�+��h�*����K@��T���rL�]�Ӥc�iz*�iz���r�ҩ
6��Jб��sU/�>x?����\;t��ʌ�4�p��g|��l*���Wo��ӈJ��$--ˇ�"�@j�kM����W��1_8n�'Jz0Dc�Hh��d���VV��Ƥ����ɯ���uUt�V�qڮv�:��pg��u�]�P���ض\e0+\b����<D��4'u~��~u���"���(1}�մ'��˫��~��g��XB��;/�UB�y��f,/��Ï�7Q	�{��� J�t�@�Jec�|xX��aLg<|�ǪU�_�UfA�D>0U��b�!q~��ԫ���t=m�����S@$�Y��#V]�Q���-L6"��-8#W?]�/S}]H��~ؽ�Q6�޿(�d[@�F�M��s�	r�z��z���{��{�:�RJ���~t��n�y��yS��(���2��`#��[�j�`���aH<�J}Ļӛ�NS��
{2�r�>��+�W>(rCR}	� <.�C�Yv;ϝ����Ǩ�ZJE�b��R�EX�Vؑ�-������;�z����ɣ��#�|}�RD��ÖΜ��⺗�F<���e��@����̰C:��iZ�u��h77�u�z8p���W4PaA��R8+�cR�X�`�Ð bQ�RYR,�J[ҾÔ�P5 ʕ��<��_I�c�� jrhT��'�o4v�W���[cⷕ����i{փ�d���E���1*�t@v-^tv��E�Uz.�[.��>̒���ٰ#�w} �DRq#"o��(����s���ݳ6�s�!`�=��%�v'E�U�gi�3����Kܯ͒�^&B�Dw,G�V6�'��ľ�ދ�BQ�.���FWR��v3t����� l}�7<\���-d)�����n����#'c-$�m:�����KIS~g[�QrN���m7'�7����;9
@c%!b�'Qp��AJ�����qQ��
��p�m$��s�l	� g�;0�x����Yܱ�ǌ�M��Q/�Ou �sg7�)'��<�����!���A�[�V}9���%*{t�YޞͿ�d��)��uGݹhp�[/�,$��o�,H���ލ�ǑU�M��)��鴣�}�vʢ5Uk�Ij��}�)Q��W��\�ר������l��gF~�
��=�x�K��K��&�ɴV�F�~�%��ų�xg%<�tO�Փ�4�����C��8g�⳹���*iϒ�ؤ���M���l-�D2�H;��w*���.7�Y�B��i�*W���R��e���������JɳW�=U��0G��Hɼ�w������dSjj�-��1�P�{�<�M�h4r%;ea�{���K�5�
���<t� ����7�N�����+Ѫ?��U�2�1Q�u���=��4k,�|�X�բ�D��	��^sM7��R�%�C% �b�L�=Ymiu�&�r͕ZH�}��?��$�򧂧��x�6�*��T��ym�6P��,д�U�����3���{�e�B�??k�Kl����g91�����]��9v���j>�>s/�JW�0�1xf5U�*dw�D�?��Ր�XLBMWǞH$��[�;���ؑA6|��8�`��r���-��Zphg|R3��+N	ʄ�����䲉��JT7��� ��XpϜ�J.*(�UI���*��E�l"�����s0 &&,1�e<�$�@d�Mw��j��Q��;'��抹�c��^lh2�$P��Vf�E�F���T�)v�A��xM��M�-R!V���-���',��缼��
�+^ٖ_�gaB9�P^�a�(�G%��k�>Xy+�*~m	��x��k�R���ڴP����Rgv���|`�rnUk�Z!]BX���u�̹�N���/����Jt ����������/�B�i�8�����%�~���X��<~�3=]�N��*9��VC�E�])vc@H�[g�ϝx-�y?�@�\���,r	`(%�m/�9���%��@Y՝����3��@y$m�?;���GnC$�o�=�h6�C/D4ޜ�\�ʨ?u*���N(?�������Y.ݿ�����I��O��<�(�{Rr��@����?ä*�^�������3��4M�C��'��X��΅�����-�?j�۶r/j^������F�.�O��L,�D4�v�������
�`�c����TF�נo��l�R��fKW�������@H,�f��;(r:������d�V��?R����h[��f�Ñ�݈��
A?Y��]�2���6>R�v��h{�1�q�7Ot�jR�s����U�3��ܕJ��-95 9n�d�Ѡц��ĞB�G0��/>�zBq�#���q��$��7�=|��Zդ�ͼ�y$`�1�Ҽ8[8����F��ɭ��{z8�i:N2bɡ�a�W�tj;��<,� ��z!Ԕw�FZo�"�ؐ��1�a��;�O���rK� �ri��7���1��K�<<�*����N�-���Jް��c�m{@�ʸ��`���՛�����-Hz�M
�JĮ~>�b?���x�[��(@;��'��7�I��H72]D�$��v��<̒���{Ϩ&�n]���D�D)R�$�t!t�*��ރ��ޔ�w�.]J�ҋ��;�^�~���~�8?�w�xǻ��qe�WF�}�5�u�9ל���L`!Y����A=O�f��0��G� �e��w
���^L�����:6rp������GJȃA�gY����>����zD�5���бXh�0l'0q �b����M+�ě����U���)w�z�S���p�r@�Kd��B�u�Ld�?���\%W>���2�*lʫ}sM�|����,��sT,Ќ����&(��%]��1��S�m�<VY^agY�l��G,'nS��4)�*l��;��=+�"�/|0�):����h]p�m��<_�O�z��ː��U��o^� Z�-m���`��h� k2EN���� ݕ~��^��_߉��
}ؑ���%3߫޳@�	�w�6
���4*\�ȞR�����Z�˺mtf�T4����ǋ���bncy�m����*<{l�CI�r�J	��B�'����� �!�݃0��)����2	�l�5���޴J	��R-�[��2o � ��众��T�c� F�)d��!ڄwJ�E��qgc���I@�*?}AV�1&SW*vH%n
vtJ�r�`���������+�y7�H�=4��Wp�hŦ�Q�~T>@r:�5��[?R~�tq��Xđ	H�`!��*�>]���f���07�M\��N~Q���ȸ��-��)�r���>��
#�����sZ�̞�~�b����d�g���>�v�r���X�F���3����qc0�ڬ�HL�w�V���z�[��kA�5NZ�
��Ѿts�u?:��#�!Ϲl�}">��{�K��Љ��L�«���+B�+�L�	@�<�Pth4�s#Ey�$�	��cw�#nw�,� �Ҍ`��fܖ
N�M��=�1(l� �z&ɓ[q�0뒁�$���u��Px�rOe���e�)T(2��F4�,��:�(�s=\������S-_�nڣ:�	A>Ch���Z]��z5�n�11���J%��7��e�Ьe#�O!�S4�􌮴ܞ�P�#�8��!)�쵆r\���9�ᨍ��5ܹ���t"�xe�*�@z��C����Č߅<o	���]�t��Gy����H=�\���V���עu�I����ٲ��\�)�EzC��W\����W��ZfI�Jf�I�r��x:�Ly�F�__r��{u}z�-:`�[Jܑltb��|�u����]�J��W�ݗV���`���O?�f$���s�*�jw4�W�D�<6K������w�p2m�eH�fbճT׼!���}^����\ie��ܻ�gS������nT.�ɞ69݅���{Xz��V��G�ל����~���DkSП�^��q��@"�7��IA괒�͕��L�W$G��<^�����_c(�E��3�p�&?~?�ȡ������-���	��3�~�?�����L�,���G<Paʪ�E�5��Sv��C�[�&��_�#Χ��r�����0{�rC����w�u��ݖ�Q���wؤ�EoJH$\i�z�Ӟ����K:�z+����%A�aod�t�k���5LpU�&���A��A��{F�lU���'v1Q�ԇ���4�(�U����뿤l�
1�bEں���3�V�Lo��!�}�7f���}�H�]�vE�q�z#�%`):Io���ͳ��$��Jp�5{��8?H]�~�gR��i!�9�z��F�J�=��u�S�ؘ�Pq~�DFP��	�0�.@f"\�}�C�!�n�
��E��fvn��zg'H�/�w ���B`��V�a�/�ȵT�S�����M������fV��	ôqL����o�gG�#M�@,x|g)��0C���?l�R���!z�v�eF�[�*o�B�>��~}\s��q� ��~*�W6��i����btMѤ�bT�rԿ�������A��a/���t�J��B��4 �y�g6dz[����-X�`}Pz~>��[������JR� �L���RZ�H��'��\D����s��+�r��c[��o�(/)[�6ǜ���D��X�.��Ő@gl�+-V����S$z�Y�Ƿ�t_�a�0Ī�����㝩�(���,����G�[_���mg}Y3NJ��3���(/�WE�����Ў�Ώ�
Ч�}��̵�+O�)�m9���V�7�Z���L��]p��Hv�3�B\6JG,v���l����yp}���$T����3��?j��IAT'X���s��<��*Vj��	�D"W��B���~I���<0@7*��!�voӬ[���ZI���q ������PjE/x��a�:՚�P�LxNS3����g��fM	��6=�ɞ�"�G�C�?sC��Ľ�H�]��b�D,�VJCo��9n���ԅj��Sn���ʌ$��X#�*�t��e����]|K��<��q�z���=/:��o9��u���-���k��N(MXc��w�0c��S�f2�p�S�����fz�XR�lK�?^��7o��t��X�U�����Ν���J�;q/ϻ-�@�J��"W�Xw�l0��!9����Kz�Jz���ױ�d	��
}�;9>�"��d�q	��ȧ��l�G�q�-��@�����GcԽ�3�~Xl[�f�+�l�b���j}k����U��ʄ�p��ԕ�@��<���HFJ�����Sfp��!?��m�!��ր)
�� X�ߘ�N���|�ҋr���T�n֜�����������/@�հ@>�Q��Hv�`��]ohWm����ՂM�����j�1�Qa�Zķ��tj!}z�'�4l�� .�#��FR2�])�Q?5A�?\���Ɛ�S29j	��Fq�̴F�+5s��zT`B?
L���/Ez�b�S�##�LǘSo��X'y�b��xPDc��5:��$�(B�Q�/,�.ބj�O\/`�|�d�j�^�ޏ���ϔJox=p������ȅ�^������T�J"����Kn�u5DV|�y�?��������ӕ����먑1<��;�,^���������y����ĒkL��i��I
ȃ�r���Z�9���*hkI�X�9���,~�n�f�
	s���K�w ��ɴ3�zQ]X(���X�3�+}dͥ��!�����KpXa�����DQ|��b�ݒ�jM�h� E��5�������`"���Ǜ��B@��+��9��O^�k���x"���4�^
��j@�I.T����g��-K�uό���z3��s>$�觐\$h�`�o��"L�VE�W�$���z�3uf�9�v�-F�86���*S�K5� G�[��\�rc$��)
'��|j(&��<"�nQ��a��:h^M�#xaN)vK�d�ٙKx8ACꮔo��iL��"���Zdil��^C�Kfkɑ*M��m�ۑ.1���Oٻ���5�����"��n�)��c%���SM]�U
p��o���C�M[0��`�)�1���#P8��Ъ�>X^g̛u�啃��F�a}�i������<;�6�M`�U8��\x
������)Hⴝ~�y��f>hmoT���HS
)�{�*�B��D�7�|�9W],�|O�)�������Z��;���/�N/FGa� ����ޫEl����x�<���%k�(�������qU�>YN�9�{��5�mk��sH2V�)�2�e�ӧ��lQ�3f�Xc�.Ԟ=���g��o;��XE`���)�d��5Ɩ��?t�oI,i�5Ys�ŗ���D�l�쏫������	W߼|/mN���]5����������FVz,[�gʫ�i ����>�Yn-�
Yb�����~`��]іJ�.�p2g�AK.�'t��J�� ]k�M-�6V�-oN���=�k���E��WGb��ʰ�ɻ$uğE� �kD;R�2�U��i ϓ!iG�?S��X�|�S�J�D�dy]�hR�h[���;���'���ز1�a/�?�tx��c$��W㆔j��%��A���q�q�ꮂO<��A�H�����a��#�O�$�$�Y�;�A�t�{;�صE��gbA���Z#%1�
=��K���S�M�"z#���W��\'0��D3�Lh���.7)h���>��>�r?:�p��c@���,���Wh�Zo��~r���Wsz���n|G2��d���!��(Y�sޏ�>����g�/vD�s��=�q���:M��v�"/����;dc����K#:ZP�ֳ���֕n��3B
 m�{��a�6IF��`T��!1{Sp�>[x��+�����C�/43����t�9��_X|޷4Tb���l���J���GR��p2�^qiц\�̂�T�jM�݆V�o흽o��y%���G�t:��)ܚ�����r�0-���X�}��=}�� B�j�9w�_��4|�C+%���$�u���f|=l:����D��W(�~8�VIj��V��
�`��@�"_�� ���g�4�)�!r�9����D��9�e�v��0����ީ�o"k���H�����5�e,���w��Ύ��W1��'7�W1�$��\�m�m�G����k~���d�80l��\�:K봮{����=�����w9��V](�
u��9����`y?~@7��F�o�+s쳣E�Y<	���b��#`ȐnrJ��kr[�c�w��ke���g��tTv��o�`�����k������l()�������`��7<^��ai+��K����B��R���_X�_o��;�>�w�ykO^���N�A�K�r���Nw��o/Zz"J��2�����r�/����`��^@E�$T�����̑�F�)��q���c4��B���.�\7��i���ؗ	�A�g>�p�KaK�ȄF�����A�y<�Į��H����<=V�g>S:�f���jm	Cm�6�n�!�}�fj���g���|�sB�H5��ל#�_�/���0Q$�#�y��c����O����O�c��0+��% ���D&��ũ���P~ImR뛡��RҮ�շ�M�٪��grfj2�2����9�q*L�Ãq���_U��3�	��&.���E]�{��IO�\ea��hԮ�n ��-�XO���
��j���vx��L�Kt��b��;M��]����xU|��tP��bUӎ���@��r9�
~�t�d/ ���B�����թ��W
�8��ni�n����F&�+��ͯ���U�&-���3����ȁ�\fM _��o)�U��d��V?�7����#w���/kY�t��zU������M��U���X�����������~@���������?E�ɡ��h!�����}�&�H�0�&��;Ф�@4u����aS����Z;h.Y��5�A8;��O$G�y:�Vr�y9��,�iͼ,Z�#���^-��݉���V�R�����X�7���ԉ��|��^�׌����e�M@�>�FҢ�5��T�����p��S�B��N���EG�E�!zY�%>��Gr�R��pr"0sj����F�L������z��P q���٬���D�ע[�ɯ��ӱ������1�b&��_8;E��^�ft� ON�X��ľ�9�L�yt��x�{-0f�ϯx�Sb�`)���Y�����+F��Z������-�s;�Y�*��䩀Vyl6ocZ��W��*�J5q��8�M8�[�X���~�BT塞�YhLi��	�/�&�:�,kygyS�p<@����\w:������_��9���Td�Y��l��l��σ�=��M�N����	��I�a�D���y�/����-�#��B]0�e�9)N�b�΃����d����sL���`������ح�[Ib��� �����<�F2���'Ka��ɢ�il0�<�[��kP���������!�r>/��މ��`�6Z"�uE.e�!w��89ʳ��p������ȋS���*�ؕ��׃��n��f��̧@��S�$��S�[� �Њ0��-^i�����_?�NIg���_Ad�A{�o g�6�fYև
�}45�*b?nA�4�\~��L�֡���\	���)��\�A�9\���.���Z=1Ny�d"�@�N/�l?B#N��%-V2��<v�t����=ӆ���l�|�� #�~3Y�i��L�3�0�W�]�o�~p��>f�SZĞ4SCr�F֮YpZ�"��ݔ��/�Kي�?2b	(*堰j~����ֻ�t�������?]ԜWhi{ݽ�^�1��>�x������%�)/�����W�z�����������4~-.ru�A�9�e����5�(�Nyo�#�{Jk�����Bqg@��A��(�~��1QI��`f^��8��"�����'���F�띦�7��]|�И��|�f����"�ѿMph���Y�`��7�����j��0�~&����ڬqI�����֗҄��U��ɳ55uO1eaVz�-T3,�"��$�m"�d�&|��S�ӤK�CD�3]�G}�A�#52{��1�:n�vM~^C:}�N�n*��IQ͗ge�r:�`����U����ke�ߧ��!Z�s�P)�]�	�j�F�8�o!�F�H�L n�Exn'_	�<)q��bZ�2NO��/\�IB�$��rr�[�&R�q�hG�$s0�����hhX��O��?��5�d����S��9v����A�O�!�mE��0U��V��h{�>׈���˽�_5�j$����x��ם�z��-hv
)]�ڃi�����@�X�ڢ�O	�!�?�̳l3�����{a�zi�?a.~�����VP���i=�#sa��RTS���8�֕��i��g�rmN�Iћ݁�{��NE��I�u�n��GYV��P�H���L�SV�Y�:�$*�|��<���q�0e�˒XL�����`Z8�����\P��8��(б�Vv0҈囼ą᭸YU�|�'�F��iư�ʎ
�h1�ŲPZRU@�E��xW{��(���s��B�4�Y�}�Gc��N0Cۤwh�D��:�����T-[��ѭ�'���U��E� �Ίư+�@��ڳQ�g$�Y{B��Ѓ�!kv����������H�'8"~#_�N���t�&2�K��~�/�ʁ�єD�^>$mu�,n�I�33W+�!��nS'B�x=� ���ϒ��3�o"G��K�w����GRc���#�#�1Kƕ��S���L﯃e���V���FM�B[��zg��`�iP;֕C��B��0��_���/�S��D�/Ǥ���mH�+���b	�K�*�2����"���`�}�!a�)NМ����&��&/�������~��7B9���ҩF���+�IE��μ9����~��o�$���N5m�w�6i��Z��qw>��y�r�R�3�eH�� -���c9X몊L��u�x16Րy�#Mf(�CM�֞q�U�����{�$�"�M7V�$��zpt�5�ǨJ�zm���xzD���z�G3I�����]����9)�Y���I���k�j�2;��I*�?H�p�冬�����Z�]y�^YZ�H+Gj���wm!4��
���+����$�ҐT�	/����Y�9���}��>�r���B}�/��dÆ*����(0MNVY�!�t��%��R��ONL���b�ELj�9���{�ź>�P&e��B�b�}X1ߞr\�9�w�s�O��G���1�?�j��1c��`�$ =���B^����}q���'��B==��P:,6Aց�i�T5�q[�����`�?�P�h�=]/��%}�I�13ݸ��A;R���'TT��ƴ��o&޼3�|l�7$3�E?(n�޼�	���ˢ��_�+�/���<�p��1hM�wXkw�2�b�����7���О�O�&ST�Bo�����^�u�����Ǳ�p g!�����r�-ir�ه�yb*ad���q����h�����|���itoJ]�H:��&��ǜg��_ש��1a1��Eq$s���|�����$�8�U��g�G�(�ܱ�Ȫ8ye���2�Fͥ�9��j�P��ʩ�:�q�&Տ�Y�R��e�=ޞ=*�}P����#��#�A�#��������6JG��l7{�ǫ3���u�b�6��炝>Ьte9vMn>��^�7e��Wz�W�`�c�XY��^Ҋ]>뉆�1�u�L��Zr�^�߿����ӝ�BG��uA/�s�:D�/k�f��%�M����Sn'��������/Z����1ym�	~����s��e:�Ƽړpp�r���r�i������jj��Z���E���d4g�
jR-��~�"V��X(���=KnH�N�Q���UJ֚�}mGaU�V(���|;p�H�in=��ъh!���j.�vk��w^Ui��#v��G��Uy��C�I
#Vn ������&$";Be��>'��L�1��^����S�;�N%��Y""I��_�����X~���虀��wg�Oр�����U�+���-��W��sF��@P���N߼B���p��쟫�4�JPS[�4��{�ɉ@"f��O�cD���I��w֔c]:�j���e�,~z' W��ݏ�?���-ִ%�V��T4U������U���xDΆ�hPs<<#���&n��<~�Dz�0Ț<�Kf=�7Z��}R�?�/�C�D��u�`	�d�P��_�B�(��\w�j�^���Cs�Q7���OG�h���V5�����ĳ��h>�-�k�����gy���%8ԧ���M�31��5��D����'Y������}w��0� ���Bw��SoC�÷�j�(R�z�M��"{2�����p��7����MLK���s>��4������aQ�o�ݙ�Z �r6�a
�o )�Y�/�v���z��B>��.W�1�e�,~3lt�c�y"�`�.
�=X�9�͠;\{QW�����oģh/�'�{g�Į#�c�	u���&j�42Ԟ��]�=.�]de�W�32�hעv���4�6��2���L��F�rǜ빁�yP����� ���$qDw}c=3��{��%f���oWso�|����")���Pz�oq��p�*��Q���ގfĉ�8��g�o�}��C>�SK��V���Х�5��>�T��X8.<Nѳzf��Y�A
�gM��#2�b"�(�+h�}�*�p��OiF�tFN��Q��@�BqL�$��W�Z��-�D�5�X�/۬OV�/��k�x���(<�m)����l���;n��e����ߑ Ur����K|3�q!� ���4��a3�uM�ꎾլ�z���a��/��3�[��ʙM���F�_ٻ]�C�-����Ԇ!�|���Lm��}Y虅�wW���@\����vW�,i���xQ3#�����u�t6F��9����j�<*��ݘwGVd�A�>
[/<���
�zS�; ���9Ec63��
u�e@g6�7mO��\�M:���Lt��UO���.e���>z��7��18S�"��D�X�4�� �'R��#j��s�����F�	l��G��"���Lģj�J�6� ��I0��}~i:5#�>�O��%�������`R��4n��{h�:�\do+��U1�G��Vm���$�KʡS�k�|}�'�<ϐb����?�u��\����3�)�2-��L=�ϒǨ��k�Y~�=R,x���SlXS��)_��󵊙�=��F2���Ғ�6X���x>V�	���<���ۦ�b�k�b�t`3�!���X*5/'(jAf�GI�1��|M_����V�Ƕ��T�C}����P��?徖aAl�vЭ��V"�^�K�f:LD�̗.�{2ڀ��j���Kk��%�
D��������qO�z����$Bt�̦6�^��^x�@����	�������`�����"�a�y�w��d���^׫��\��x�#Dx���Ʊ����V(h@�Wۦ%�E��{q7��k	���8;Mo<A S�9�՞�9����r���UD]��$'�3<";��)��g����L�o C���3�
d���;�3ܧ1�)��k*�9�o^R�㽨G�g�fS�	P%;fX��w��y6���3<k����p�[�Hw��+�� �W)�V��JL&�(�p��Ƞ2�-@$2\��`Z�w�z�hQ���BZ�~��v��Ly�8&zbMt1�vP��TMM����?__�EJ�t-)���7� �� �UUp�qOk���X�4 �F�v�Z=��~~������b�h���hF�s��o�tT�C0P��3YǦ�V�޲��Ж���VV��K�����H���G���B�z�Th+�O&�����E��]S����$_Rz�ʌ��Ǩ^>��|9�z&d�u��w�����|L@�]Xg�X|@�x�F���x�"��Ƥq5Ҥe1[Gyd�d�@�?����+2�������kDMv�h� hOR�Z�Ӑ�+��%.��w�uf�d�ɽ�bp!3>^��������<�!�b�9 E��ɳJFa/L,��`&��k\{~����7��;���i�]�2�����$�k)����w<�A�9X�ߗ�����A�ka�2���7�u\��̮��e]wmS{
/^�}u01I����~E�m�8T��V�ޮ\��7�ה��2��� ��z@�V��.�L%T���zm�l������$s�1��'�}���y�\a�b�;��Ɉ~��';���I��c�V���gJ-WYk��C���L BÁ�'�N�Z��KnK�T�	���� ��Z�����L�N����VHg���lYV�Ҹ��8����	���yA3����4����h���Gd�<)ey)­���4���ɰ�t��$��Y� �F���m�`�2���!�+��=3�1ee�<b�=�I��gW~�&��}����!v1)��L�[�KiZr$��ڰc�8\Q���0�ZwbASy;�̅�F���B�z�/"#��uj�v	�y��2xW�%��K]�6P���ֳ��^��c�2x��幅�5<��iB�y-���=�V/��J ꮐ8�2G#�1PƗ�)�b���Y+�� ڞ���-��4h�������#�p�Gg�,0���BJoh".�k�}��t�H��%�)c$m���n�����`W���Tw�ݎ�ю[�P5I�����&�'�x�"��a�-�����ȷ��tѦ�1�;�i��4�,�W�_H4��#�C�[�ɟg|9		�d-p4/�p�h5
�8���~\�R#�4}`	@6�Խw,,���������=�P�ִ�v��G�=��̏[ѥ�,f��m?�e�}6�v�>@A�<��;�]#�3�2���¤��%)Ke~�yzY��6 ��;}��<����C8h�o"�a��z���	p�}�$���_�?f��z�=<�f/+,=��?�ƍ2FWȓ�������~Wm��Ϥ�;C�6/v�T�Ai��B)��@�w�U�\����Ȑ��?^��!�]4�I5�oc��_YȂLߏ?�O6�}1��򤶘����/T�����6ls��v�g�K/k��R��O��*�I% D�$*3I��V=��ܫH��E9e��[�9U����*`c��L�8�kq�94��{����Q���B�����c`�F/"��)��=PXfp�uC`U+��:?���;�_���u\���]?���'�r�H�����ߗ�C�嗏r�p�+�����Qo�f�:ȧ�%q��A
357/LTg����d1�6��8ݭ�����؅<[���R�~��/�]UɽC	�ބe��ЎZy=~�|��W�Va$����&��"�ö£�3���1���q�d1/�z}Y�^�H����^Q�K����R��o�H˳�u\�Q��AZwf޵�(K���9��J|�_�<�,�h�V:�D%[�"lvU�@�/B�y����v�v}9&;�e��"��`�!=��q��� >��:C*sP�Tti�@r:�^��k۰o���#/y"���.sT���X#�0��r��Y��H�0���a������ᇕs�C?[�.t��x\7ϳ�jD�	�3D��{�o ��ꁌ8Z��{/���I9$�yP���DBF���B�F�#�ȣN�nw��c����ޖ=FG�P'�v=����P��n��ױ�v��O�E�!�DnDԃ�W��>�+ݟ>�w�(}P3�_��|ZKd�7�l;���ݡ��a��J��ܟ·j��p�tE����� -�>�j����_�Ц�yԑ�v3�2�*�>����˔���/�<D���fa�c���Z��v������<ة�dGx��e�Cfb8�'K���#%��xE^�c]4�QJ�}��å|K�-��aK�`������8q�1�z@;��vņ)����"�5������5��^�o�U�-w\�ĹQ��Y�M�,p�,���Jk�E����.�����tm�$�X���x>�%�����~�w�^���RM3���A�\����6N���1�D����uY���.�?��/�_	������_��'rEL<�P��	xn�d?��Epn� ���V�������$/���d7 �I��:����>����)������4/��P�'�%�B���w�e��Q}X�Ç�oKE�	��B`�H�b�5��� qz��AAl�!�Yձ�|T�_�w�+�^M(�5M�g"Kz��`�B(����̟���0�ָ�m��B��:i���&G�9�ȭ�%Z?�F&yz�#+m���$]h�Ш�D����!Ǥ|���V
;*���ݍKU[Oc�|4��&Y��k�ÄҊ�KSp��q�#{��G۲��#D��&�Mfj�av�Z[��r^�?�~�e�[p��I�m�G!�滑�	�]^�㉻�-��F�����,
1mH�Uu�G�uF��zV�W��������R��NJ��|���j���3\)f�DE��:�&nމ�{����E�������T,��t���1�����pn�OlYg�.K�L��w[�P�t�C��9s-\��>�Q�3v�ۄ���1nv���·d.�ӶP_�Y��ۤ��Den�����~�H�[���}=|Iy�5\���	Q��2�t��g�W�k0���Z��
�&����`��1�\�Ut������U�j��R�LW���Ki<�p3�^��}��o�n|�i�6e!*���7������NGp�.4���-6�?ږy�"�9���F~Awgţc��r\�X��� t_��|�vہ旐��H ��u����*.�<;~�|�����]�Ko�����w�&rޏK�����Qbj�#y.u��ߡ��[p�Ax���w^Q\LQ*��Z��d�}�[�Q���`ɛ���V=+�:۱��E�M�V`vn��0$s-��kZe�R��͇Nx/^E�Nn �6�fa��o�o�������8��'^�5kӿWm��;�G�0��?'��1�/Ӻ��W7�v<q�.�ptBA��fLTV��p�dSm�G�E!� ��MN�q�,�RcЗ	����F���n���Ű0G8�&��b�p�x��/����G�r�5f݊��o�=�z�k�
��]���a���Bc=�K�d��d?<dH-��ݱ�ۻ*�Ù����^�k2��{%Y��ƷTq��"p�D,x�<���̇v�} H��ղ��5�=h���E�R�_ǭ0����a�WG#D�����7���橿�ۦ����L��ih*�:E��n5�0��&�G����!aV����>o�T0g�_>�<�L^�1yD�hZK�n�
�75d:V���r���`0���ǅ�Ĝ<<�"�d�rK�1�TL\
7�~�+E�=|��B�T
��˃����אO�=�Ռ�vV�t�B<�"�ԇKOHW��٠�{?��6�GlBso�kEs��ؖJ�c��Y���Ndty�MQ�m<���-�4���;��+��C$_���c���h�s�
�p�`� � }/�odLo�N�)��/ּ�	��|�B�E��q����G����L}�����D��3��v�ą��C]����¨���,Զޡ3�N��%r��Q�}x��E���e�.�y��ʌA��#�i�rS��K�}��L-��Fʇ�4[j`�ߚ�Ƙ_����+9�Q���t�ۮ���pN�8��aI�0\�H��	��W㘛��������;W����o����A�b��UAY��x�q�>�����4Iw�E޽��&b.{�͜���n�1֯ֆf��#�<�$H�����%y��e�y�࠶��D�Y�g�~S���g��WiG
9�0�co~���vw�����5j��d��7s�7�Tyb��7�??�/����<����e��*-�(D&��ܕ��1P��@X�S��KG�jo˗��'�qRx��CIt<��Kq�/v�������0��:y_΄\��$���+\���XU(��~��\��ku�x�+f��'�[K��v�s{����_�h���'�V��©����(��>�QNie����<R�v*���y��!�z[UR/�<r����z3[�[:��9��P�z��`�Qߛ��'u�O�����E�r5�}��XhQF�oU����5���%��	�c)�+���N,QQ�d��2�[G�B�=���e�l�.F�Yѧa�*��j꥖M�D|���ъ��X�a�n����J�$`[l����+�w�:��s�%���S06����O���bT����yZ��W,N�,z���`Mo^�݅�n���R��\qWx�n��������:�D)��*)�GS�p�C�����C
�q'�7�Ӟ�wK5}ԛi����>]���k�ñ��\��{f�@Bm��G�e���,�<ie%�C���W�8�(�	�U-44wu]&�'��1�V';���������Js�b����4��{Z
�Ƒ������ܳx��n�^ί�o� �����k�7͕'�d���6'X�R�eԷ��d�;1h]D�T�����d�1z�s�"�)h?�m![�V��w���r;X�"c�E��yD�u2Xp�(�n�a;��WI7du=�#J,�jYկ��4�H��Tn�� �W�u����Ů��Z�Q���t<(�u�P72S!C�4�c^<.��cFR��B[� �Sz�k�K��6h��\�(��ª]��/x_9/�'��2��R¿`
w4�!G�L�����j4����M��{���Ǆp�t�f�z��b�J� c�>q�;�tsuM��5�oA<�35��;�l��ѯ��ӄ�����B9"�������Ä@�߲u/�?�!�lw�\M���IKK�li��ST�� 0���D��i �q�U3�ٽŋ�6�i;8�5#����s�*O�v�ZW�Gzo�s-��|c�w�����M���k�>�̯$�oV�lQ���ǻ]�?;	�>�<��ń�e��R^��C4��*���p�I��$�n _@Ly�-FxpFp��nW�ۻR���Ɵ����������Y\�R��wcB�띜?^���lFK�ܭ͈|63�&7�n=$w�$����}�.��4S5ڣ�k!e
��W]�� �oX]�!�aa��6_� �r�;4�^�k����G�A�^��������?%���a?��Һ���h�����$EQ�?X����!��{C�vECz6��o�l:�d�J�7�	4B�[ ����TK��va-�(|#���s8�)�$�s��Ԇ�tt���2�7�.�R��^(��l�kv'���9߿7+��625) &�Cx��U+MU[�r���T���eU��T8��`�8���id�N�)�;��K#��\��Nr',����x�:��½��қYV�r�޴P�/�]Roe�BS��=:�k�a0��m%ր:�k�ҔH�Ӯ!b�~ef7���(�.Z���%k�j_�'��D��	x<�̟�=��G��C��M����6�LL?o��/�9�2PԆ��T��?����C@̝��!.�	=Z�Dw\���,&P:3�.��'�<��/��<}Ad|��B)����d�@�{[W�Q9�����	Y��Y~^�W�ޅ�q����]bb���ߵ����B�P�E��6�����X0�s8�(��(���vFL�Y�%U���s����߀l��~3�ô���F�7���G��7�Ҡdh��/��M��gS�B��&�v�Y�����j��d�R��a�͟��>�HnЬ0���PL�Aaw*�	�|e�w�N^��G�T��z>����6nl�Ov�}`
���	2��6��U=�z9�<Я����II_�hAr���]Cw,L�O��~��(�gV<Q����%8��T�ד�!���� <9�{�� ��>H���b!�b�����=�t�m��d���� ٲ��)@T.�^=d��޿�_��'�x��JF�`�b�\!^ �O<�l�x������I�=��L��CO%��9���4��V:Ǒs���ELI��J!�y��Ψ;���8-Ĝ(�p�z�w+��v���龏�_�c1�B��(C����!.1�C9�f9��0L]9�X�C1��X94"wZ�̄-g2��lܮ�q�������}���/x�?����>|v@��L�������a���6$�
�Y�jY,^NVg����3艏��!!Sm|�v�<�8� �'��mH4U���:�-��y��P#_���v��"���rN�"�q������,D���z��#�~��^��7��庘o� ��J��l_o)w���G��"��K�S�qY�\U��S��!����}#8ߦݜ~���Y��^ӗCd?�3�WDz�}YJ�'^Tf��MZ8����
C��.����?H�W�FJ�%�[\p �6R4 r��r�h�}����Ro�=���,`)lW����c,�@���С�t��E��V,\��7N=�J��.)�#�G�Ϻ�t[�|fԘ �_�$
{�B��5-"!�c��'Jw����;+��M�Q�.�f��˖��A<��,��&d�0<5�<��\xZjW>�@Ok���΄����#>�8O�)���w�Q����u�z��F�7G�����v�G4�����ݵ����vrr9sa�H6�ЂX�2�4����HQ���~;�� "8���S�Zk���I��b�
��P|T�i�E�"e�6���t��|b-����Wwa�rv���<�s	�)�2�\��S��
E�9��ج�w�"r�&X'�>`��H�e�f�tw����:���o__��~>:�F���k��`���n����%SC[�ĉ&'��2Ã�Ҍ�k��ޝ{v�qsbj�ox����1]������hYX`���l(%�i�<#s/����_P8�Hc��Y�{�w�Չ��z��ՙ��$Y7�=��3�����N�	5���8i#�Yb�ұ�ѧ��Ps��k뮃�;}�9�EWR��o\�]�ASh�*"�/:Hm����������w���$�8�˦�'W�xj���VYe�K�(�c��
���+�"]xVN�gFc�������BrB�}"���M	n>�,��	v�Uj����R�؞�����-��cylk%Q��.�c:p���+��D�Wx+�P[��� ���*wS�'��4����cw��@�cp��D�io+�����1Us��{�����%1f���s�\��xF�&���|�=�p0���
2&i�p�����)�㕼Q௑�ј�2����]5X�lG5)N�����Dn����e��}:ߕ�����ƭM��E^ P~�M��������RQQ-(���8I�Q ���9��NJT�M�n�8�� ������̎�;@_xz����T�8�ū�]�}|��9!&[�u�Yvŷ��ZG����!�Z�X����Ϡ���'=��*�x�xF��	bLpTӒ�L��Al�V�*�d88�l��E��<�������|.����ń-9)�OIڍTR�E]j��%��3^'����s�;�j�*!	C�Ӈ���3�؏�Bs	���<=:Ì�R�0��{�bi������Co<�x����3��FB �u���[�%�u��TzE�_	KSA=��>��d���=⃈X���Ȕa�:a�X,G+�LxgY��ع �X��*��Ύ����M*LZɒ�DOU@U�ٗ��S�v���9�S�pm��b
0b�F-7���ٵI"*T7��y�
�.2�V2�L��a vlIO��V;/����ia�8�~0��U� �4>����=Q���k��&�z� �=xԫfv�E��t�Mo�}i���~]Kl�et�2��~Ƀ���qJ0�h�X�ȋ0$��������r�/��Y�x�ev6�p��ܚ�T�q��I�Tpb��ҍJ0�DC�����f�q�P=�{�lg��?��:5���p�?Rʹ5ԗyCAS�5�eT�Q}�O����h1x+�%��$�aO=��MA%Ng�u\�(����+7u���)����&�=�X?���$�@�����J�[(������Y�g�/X�h��?��E8y��
��̹����I���Q|ʁ�H���R3�OuFKy��V���Fz���� ������t�)�>��^t�̤:���0����#�Bljw�������l�s9G�g%�IO�̞ē�.�����ܝ���D������=䝦��a���*���&�ؽ؁(>Z�=(���Ex��G��d��%�&"BոKl������>F.�|2��Oc����~��+�!�F�Kܐ�v �j_+���������2���.���	d�&�Fk
�a�o~������Տ�PK   �I�X}�� � /   images/5874d651-dcf0-4a98-b8b4-9fcbfdf83d7f.png��uTT��=�t7� !�ҍ" "�4JwwR�"�-R"��� ���!!�\����~�y�ǵX,f�9�v|�{�c���L424��TNFA��@��P�Wx\+�/DG��j(���Q0��NN��l��������I�d5�TmM�\��!�����6����v�����"d5䩌��[�n��N�kҭ��8&	?�w�����xXh�j�y�{����B3J;���Њ�4-� ;I���TJ+S�|�9���S��������P�L��2��>S_�D�Ǌ���>��l��ڟ���ڸ�*�������tq1dOɑ�Å�_�@��/�� �(��H�ER8v�):������W����W ��D���ӧ"�����E�"Dl;H0\�~����`�(��S���ʜ��*	gy����<�J�9�ڍDf
9::jqlhدv8o�}?ޡx.��r8��4�>�7�ӧ����ĺ���%�!�#�p�_F�O��?הa�e��p5�\N����o*˵�ru�av
�܊<~�$Ѧ��!���>ʈ5't";���Vd��+e�U�̛��[o�z��-~����,ٰ�ή�ᱱ��EO���<���II��ZcY���cn��t"")[�$��B��Jů��He�HeF��7
K�Zs������4����W������a���A�j�$���[�9v�����:�ܽ��)w��]+C+/�9�9���_vv8�z�����#"�N����&[�$$(>>>���0tsK��H|���� 9����v�Ņ �e�;�";
���2V�7u�����X����Û��t�{���#�ө�����~������9��U~2t�S��qer�&��m�͎���\Q$�i؜���GV�1��a�747���)�,���>Ө9y�K�a����x{��5�H�W<� �}��U��C���f�|����H�K���j4t�2zT�Q�� �ř�([���Z�d~[��xH�	����#>�94�#�ݏ�#��E`�t}�_(��[���AXVV�4D`0��X�*`hhx�w�{G4Gӛ:�W�{{"W��E����(�Fx�񀄖�B����F���2�H1'Vb*Eے�������n���_Qg�%��������������7"aSu
�6FhW��������'�Q�i��RjF��t�մ8(PUÎ�Xp]h_
�M����Ѽ{h5��0!���(�|�QØh{���̇=9Cp�Џ�U�:�8լX�"�Dǋ�/���V"�a�Ѻ�p4:�\��\������=*[&�R``�;���ڻۓ��ۃƾׯ&d"�k����\�L�[Z��+�lܲPsK�#
�B!�б���/��
ܳpѡ��g����O�9��,�ϟhy�YDT^l�&��v�1�3KJH@����=b�!�x�W��ގ8�Vv�22��ʦ�ϙ������w7������� ��}�T%����^iH��dL�p��w:	���-�0�C|�׷�=��rxt�Rо��#$,�h�2X�v�iM���8����{P˛��>��|l�`�S���۾���?~� �GY]�	V�m��� ��{�[�i��Ԑ�^E`z�FF[.��DHe;:����p|����-���'ևn"`+1w(�����|jvU��zFu�p���f�M���3�LW{���Ɓ>��HD���@b����.d�X�xv̬0p:�ap���K+9Qs�I1<�e�bw9jW�{��	7�������l�@	�"���x��MJ�Ch�b�[����alw������̒C�\c̉����ꗱ�^�A����A��1�R��3�}j..\p�23ǘ�X�}qlme$�}YC}����YF).|uqA�������f'a,��zjc���(�wO��h�k�fH���sj�Ȯ�0���]+�;`ە���#2%��\���|�\vgQ_�~{[__?J>w���~����B���v��B�M.~���G�����c���P�;ع3�F�lmm}..���2���\:��̅vLWZ�rƑ�6�XQ�͊��;^N��͙��x�60�&	r�=||��������?m9k�ˈ��n�d��dVW��z��
_	,��2��îT���&V>sb'��U�cAA�S#���%
TZ��2#�����Đk?/�_e�r�~:%���+-'����LN�y��ׇ^`^ Z�А.1���!CM;	�{׋��׷[����d �M�9�`r"w�'���tF�X���$F���8V��2����q$be��ȱ(o:8���0D���10��J��Ky�6 _]On߷� �
�����ʏG��F����	�F��
J>�i}3�YQ�Ъ�93s�4����R���Q�Z���$��0ځ��vH�'\�cx�f���ke-)�Ar�.S,�Xy'��Vw�<A�m�%��7�+�D�$�/��>��o��ڙ9GD����c����uq��� �H�>��ͮm��!8?����7ܕ�N�~��,*5��@ "�������1ۢ]x�}zH���ST%J^t��:>b�`��h�=��{চ	�磌qs[�=�6�)��F�ρ�����l�58�S�u\�T"Vo�r�D�V��a�g�S�뛛��^����rG99��^g�*+RpDࣴ�mow��g\w���֡���iiz)��S�R�8ʪ��F�`�5:::8��mq�/e��jNK��	ؤJ��r$kʆ�����x�����<�,��Ё��B�#��F�\��~����{qq�����B�lm������������f	&������> M�/3��ǮV�I��͉�� �\�1w��Gd�%D� "GD�+����.i�n/����ĸ���'v����FL�pl��\��b�2���%������9@q#{�9�F��- ��������)���K��x�Wg�_��xG��C���"������R���qG�k�X��jݖ{W;#V� �V"��466�9�����J�iۣ2uݭ�1D:]�xo�Z0M�..R�X�V���a�
ҝ��B�DI���UTZڇVZ����A'vI����#�YҀ�V�7�u_�x�����+C��~�u����ˇ0isR�E�����v��7��Wk+F.i��h����aD��%�FO˓�F�Mu�S��;�����P�2z@��� $,��i�v��D����ʅH��������5Z���g���q���܌�OJ�0_ƅ�V��qC*W%���+���ґ� D[�'Z�˽���q�{x�><�����@x_b��w�6 ((��Q*sH.��#��ox�"����k\�
	}."��ow�+퇺���++k����۳��^j/��-����M� �T�̵̿Ŧ�.�6��H$���Q@�yη,�G���d��l�2#ԽQQQ&6����w��X����^2]Cw���������zz�_���aW�T|�_�����
�n���Aa��^R��%u��rE���o�>����)�$�`,�rG����������n(�]s�v�D��ڱ�ӖKLl��28[�	U�~�LӲ��eq(
�΀X���E�Ivv���A���1=�� U��F�9*Z�n���/K��tϕ:�����5���qS Ѕ}�L#��LVA�H���z�N���Gm_�
ت?DF�,
#�_��~��(_��t������,����7-�sҘR�QF̑v�P_W����̵?�N�*���Gô�����V��s
h��\��*Qhӹ���l9�B���E��FL �#{;���`$�XegE��'�A����j5�*cq�L���iK_L�^p��J�efF���@u܀�smb�P����R����T�j��s�� �(�Q%�`�,l�o�p��(Z���G#��ko$���5���O�S/,y�����V��G�j� ������,�˗�].dc��HlqEmǓ�g��E��S��k��Z2W v{+�tj�:�'�����;���;����K�3�y�J�����s5�}��v�'e6�S��S�=��(�4�B¯�]3�g3�_H��+)����JQS	/H�=e�qt�''5����k�}�������4��"fd8s���'��i����_1����|�Nz`��I���(���r�R̋y�;�%�'O��4�uR�Cl��po�����F��v�$�I'��P��^+~i�<GO��L	��(n�J���"I�� q�w�@b�!w��қ�Q�O���ȯ�'溷]]]G�;���įj�]����c��0����F�l�-!�R���)��Y��;�sy9���c��7³l��߮c�V�8t�b7J����b�<����шCu{�������Ro������b��R�	�\޼��sR2kܳJ/�n��g�����iu�8���dvּ6�,�A�Ϫ�Z�FFFovά]:���A^Xy4(�g9��iɟ�9����͕p�I1�z7c�٘���ō��g@j���N�6��.����A�!>��X�m��P�P�p���C�ί���
ö��^��C{HjY�+�G/�)` p�(9�
>�<~3��ccF�NJz}��B�Rf��J���K��x6b n=�>����Q_��뵉R7�ت�7�nQ�Q��*��w*�@�;��J2dI�n����	����l���"��itX>� |)�Yn��}2[~xvVuU7f��sw9xy~�V�@��j� h��?	{�+)�3O.��+|x��>腖��dAp��@��_^b�=[� 6��>���v����A�	������;l�cU�g�E��/��vU\}س�<e��GqC�7�,�X���c��s&��'���K~���H��!·�=S����D!��caHC��ΐRQ=y��P�(��q�'O�Dh���v�՛]$_���{�/UE�G^p�*F�(��n�waMp���08���T�>Y��/:�FjYR�����%���z�������|�7��,+{Tǿ..$rU���pR)��Hb?��g-�����"������r���tEJ�Qg��*�G�pnb�қ�8W<S����G��	��|����.�Y?����kϑ��7����H]��.++�r�	�Q��&`ߑDi�W�a i,� hcE�T��k}�G��ܾ+�H}5��h�I�|�g�����"�G]}�����\=�g�Pxti)�<��ok}�E��ֲ�zM3�ń��b	c��ƈ��05u�U^�O̮��s�ԃ��������.$��|��b��-<櫨�����Ф\[�a��RN���P(8M �#yE�vK��c6>��(�)6�"pYr��0��m�U��tP�^;=u2㴝o`�ľ�Ùw�q�n�r�Q�����v��)M�h	�xi[�7��L7�g�	l�L>J��6$��IF�N�,س�ۿr��^�C.�W�8�I�_���q�r�T����2Y#���!#�:'7?��
�El�p��vu�E�.V*Z�v&JW�D=EvQ2Ġ��Ų��P^ϱ��ѱ��5V�:3\�5!!�tsA�k/�5����'���1d:���r6Wz��/��~�4���m�s�'ܺBBBC��Y`:'�������$Y��2&�sm`�@F;��\�����#��@�9���'�� Ƙ���د �~�s���ӕ�/7~lg~��q%�yt{�=Jb��<o�J�,-�����6�(QQ	����q��_?w�&���Gy𸙒��8EDVW���cХ��J������7�\����Qn��� ؉C�X�T/��4�J���ۭ������O�=$
+���Nq��ơ��tu��!U؜c�����g��=/ZtĲ�+;W���*i�CB���A���圼#^H�H����Q�c���J��[or���ML ˆ����*�ZIڔn�`��lfB�f�|��� ����m���B}��~�ÀAK���""�af�q��Q��[�&����mS�`́Noϡ�N��Z0&0�=�a|��`V� "l�I��6��bx�k�����R����ޤ`�f�'nל���le_���  ���n���uTjjD�>�����(V���):)���Q���^�k��@'���r`�'c"8~�� ������7�?w&H���C""_v�FE1[~�����r�^xddvݗ�}��/DÕO��U�Jq����/�u�H�����Ag��&'���h��x����f�uc�,��uYq?¼�ȶw^D��<'*MJ"��S�+'/���9""�摰��H�f���y)�����|�ڱ�;�@�e�Fޅ88���~	ǘ�P��=Ïq�;8�m�H���T�r���4JP�^f/������nb7�wi%�&"��ӑP���~��222sd���qh�33s�z���^hV1))�o^Nf��nx���iFf�C ��؂�3EE�,�,�����6\4\p��*��\�q��yl�
1qThdR{Q��,��P�y0]�K.�)"ei���'So���ϟ�lY���P?�K��-�+�k�a�k�L�eՄ׭��B�ٶ�Q�v���d����^**��������$	�&zF4��%��R��/��ڲ2.r�=����n����#U���Xl44���l�%���8�N��/&'�L-�&7�7������*���#ɐn=--2��ǝ��eo1�����dޡ���%�IP�h�;Q�ö7���)9(�>��0RԐ�w���R�ꋟ�^A�G�KӲ"Us����R�ۯj��������e�1H�'���V�u})�d����g���lhHW|�F��}	؎�t) ЍS�����rOl��]F�.����Rhb�ع�M�z������O4k��_L���1u�u-F��/�p��I�!'��>==}.��]2�&VC�F�)�mV�E��Ѽ��{��`�����h�j��
�r��)�|b�WV3G{�m���ρ�i����d@9��|�R��J�\�z�~��/�s��4h+�a�ʠ�m���9�3GU�{�Ȍ���%��HR�d�w�7ㅈ-'JR����� ]^��-�x
��L렗�[��v�*|�~�'���Y�q�|ͩ�ݩr3[� ڵ+?���$Κ�#[[[+���� ?�r!�VǑ"� �,h��� ���Zeァ���rG��.Da�M�	��. �ֵ��6�j��T
<���T�O����VVV�V~N���&
'��g�<����U�;4E��	�>.���9Pıi?�l�����L�$�"���������0'���A�b�(�`���~@dd���S<^�O�*o�pg�M�fX��t���$��h�BA��c'�Ta~��h�2]C_�ݣU-�Q5��n �'��9�}��6Y}�2�G)�����L�G����
Q4��8��'^����١P�Ĉ}P�iş�SӞ=R�k�˙\��6Ei�Œ�Z��3���Q�A��z^�зN��ݬ����:p�̲�%miT���k`�vu����'����z7���bC�x9%���F�
���>�S�*�4]�s�'b@\�L,�]����^��Dǥ��2,�t��:��u�wrq��P�#��(���@EE�Y�!&fVy�3U�A��خW��U��<�q^e(:�ي ^�2��ޓ�;?:¿����?FZhn��#��Q�O�v�J���^�i	Uv��������2��mJ&6�Zݎ-�|�޾o������𾤅�[Q�N۫X�����>�D�r?9.bj�jM�#k%��5�a�]T��ߨ�F5��[_T���*"�@�_@ ��r�j�]��&��5��]��������yd�?� wd�`(T <����Pl
�~���E�ݎ�x���J���F���J j�����_����U�=�X�� ((8���6Ez�t}R��*��5� �'�%Q��r����61���e� �G%=����yp�I(2Gs�w�B6��sm7e�^����o�,��x��_�z�C�k��j�/�;B�*��$%%��?y��ؗvw���r�.ǒ/2eFqY[K�
c�d����h@Ӽ����`�Z{z7韮R�;<H�c�P>Yv�4ޙI���r������459+���z(�����	/��}�M���^[W����kI��1=�I��L�W�h�� `e�|�����+�Ս��wU5�'YX ��\�AS���c�DEZ�/v��"7���5��7��ֺ�J�T��`�F��P��ڷ?e&��*��n�y�㘀k\?���Za$��^��������z�]#���47��	��xEu5��ԍo��<�������8C��iE�Y���F����ZYm3�K��.rs����W�$���j�DO���v�@$*3���L\�#�-��~��4G�"��wdإ������2� 33���X�ssv�Ł5�����=�ͱٻ�����E)�̓E�i�%C��}M>iP�c_7�ӠB�ש�A��+��wP�f�%RQ�682���e��n��j�jl__�0us�� wxPm��!���&�ӽ�An������;NO+� J�zN[����w���D�vq�v�������ވ����r��3%�����t���i����y#I�/�q�������ʝ�	S�	�|hh��N�h��Ѳ,y��ɣ��pӯ$&M-*5܂VjD?P	�����J�/�K����������$pt����1_�e�N�;���sWS�k�5�R���!���
�og 
�w(v����x/1���{����3Qqsۏ�A��2�߶�GI�osK�'��
L��
��R�����%"<ܧ��Ъ���M%@�5�*���k%�ۺ����ommIJ�E `F
I���GX�O�4���<x	]�	�ry��b�fI=_��!�nC@I	��[��mԬ����R�"f��L��j����]O��?`�����3bO�N�Jx��l�8��&<�r�i�#p����0R�;��A5"@�K17�����]�P*'���H;��G� .��A��A��)�_S}ǣ'W!NB��)sK22��R(����@k���4�i��֙�В룟?eK��lJ2�(;d�PA��bѮ�[�#��V���9��)����5�j���+5�Iܕ�Ca�Ė}��c�����p��]��wP1-���c&����QP�1�@-��|d����cS�r������w���D(�Nb�<���Ͼ�мqR��Vi9�c\�����xe�)�&]��@�q�8�Jč���s��s�����[�nR �Q00r��A$42��p`�AAG�W{蜈`���@�744���/"CV���x�;�골�DDȍׄ�)D�+����9���uLK��}���1X�MD�2���e��������8
..._W즰��6dvG�>��v�(�����N�;�GP.;�/��˸�P�ڐ~,,PiNMqV&�8?~|���>�
�&��!q򘞀�}&����@��{�-�&���Ѹ��eè��� 
��܆�(~w����>�VM%B%��:��1���01�?�����{jD���|�ѨPC�Ͱ�䃬�D��>���~l}���"�\w�L��k��L$����f��b�i(jK�x|J֗2���%'#5�%�d����-�v���DX2[�~@�EL�}����n��m޾��EG�G,֎�.���:�������i:�'�cY$C\rr�j�o���Ȓ�`�T׋����{d�pU�=��&��ؽ{� �[[�R���t^A��D��C�{�������7\Rrr*H�'�_�^����Pf}Y����*���$�^~~���n�<
$4��~��o��8 z��|g����MK��G24�<-��.
�H��Ҭ�����q� Byoq�$&����8���pII���XYax��
�{��I/T/��6#4�f���gh��Q�k_�pwF���H� �{+W��H��PrM�zr��L���:�X>s�.Zu�q�`��
#dQ?=?�{�̠���{f�
X�NK�Rn:���zґZ������{"Xs��ۑ�;�33��Ƣ[���	�,�
�Y����Z�c8��D+���#��iO�Cv?@"��^�$t�掯�1�?�J�徊��FgfX�quE�"�Πz���K�j�����g+�ܧ��XH-�QO"UǺ�?������jq} Y@˝ �Tp��u����H��,��y�M5�4��7x��Ѽ� �m�T���PK~��w����<؛I.i,�+�z6�@Jj��I�o' �P��ٸ�OXũ;�Zq�4:1V>]�L�#��#iA��zt�ЭZ���ݔ&B^Y����A�+����������oYx
��c]�ӿ�&hik6J,���6 S���29�y�)~G�ŋ�����?U�{��.^e?3Q؋�cc�d���8�2��z-���b���+��V��z"n�--��x���lp�ԯomy�4��0R\)ل���=B)E��c�W>��b���xGI�(�ܘ)	�iॼ���>0H䖏��p���lgJh���r��j/_
ꭟ��9&�TT�	���H���m�e����zNM������CT����܎���i�<�������^��ZgW��
4t"V���9�S���»*,�/��!6�b����|�LF4�K�a%�"�^���!G��O��x�����\���;�(��)�+�Y׻��e1z�,��_��H���%�H�Jo i��0(=*��w�`���9����@}��~о�1���~��v�*RkO�ײV�]mw��z8D��W߼ޠ�"��apE�;ަ�Ĵ�X�7��FT��@ ��g�����	�T�ssfff2�HU�*����ֹ�d3���nPr La9/�ڦA���],|S�zH�����v��G1���I#��R�.''Ŀ�]Ϊ������h9�Z8C6a�; �Wvz�\��U�l1���m�� � &�n��Y�����������Q��:�c�[|��Yf��-�c��̃{�Qd��r�((y��Ϟ��V�W
��c�AP������������Q�}�Y*���ud[u�u���?��ؒ' y�|[��O:R@:ý�����R�tѥ��3Y&h��V�OJ�4'YK��ube�w��yy겖M;� ��mqݚ��o�V�4s[s��5�����*�f�"��[����ZOEHʟ!;K|A�X�յ��3ll���t�A��.'H�1�J˝�Q�9��<�A�6��"����V�߷o�f��Yܹ��mmm��tt����w�E_�s�sQ�(>���N8$�X"�}- y�w�ki/-��?�zN��7�])�]�{�ď�_X��� ��l�V�N�!��tq��IF��K����dS�utpwf{1�-f�`Z6f�W�Z�$��p;�Lr��|��e6���>#n���F�;�+
x_�7\,�J���L~�F8\��qؾ��q�O�O��hDD�~�"M7\�(�k���,
�׾��2�P��1ړ��`�Tb?�G��^b��on6�����Q�RS�_S�x��*���466r�Xd(w�V���R��k:/�
Y���_����=ϗ�a���	V3�2���c$Y��$��N!���aYR�������U�H��ಣEק�o$�z�G.���3W�r#�j^hNnn�v�6+�4P.[A�Fܒů3�/�y�^�#�O�M�hkh2��ږ���� [_�
$E[��9(/��5A�A~��j#�%B��d����ט-�Ĺ*������yT��/������ī�7��fhv��c[��s���ED�=}�H/��G�Z��&��^0%(,��;�ϑM�d��US�d@ڙ���g꠳���*DeV(*$�ߛ$2��K��脄U;��>BN��"{��#�������I�����H�����7u�Zd;q�t�L*j�LO��]{�b���U/ёt~I��HC)���$X1�Yĳ"{��}�G��F�H�|[���r�;�n:pPS蘗����m�&��1*7"R����o��Q5뇪��@���ǒ��P�rG���6s|ǩi�j���!@�x4����N�	�Q���� �i8;�2����g�w�+�J�k��TQ���4GC�f���6��7<�[h�����j܎h-���fHR�L�}���q��qH��#�g�D�g�2�Dt�6�J�"�;>Of�K��6��It8q ���=�K�!����UX�~�-�
�����Q)E`IY���"�0�8g(_�ɻ��+(�F���3]k
 Z��߬�M�3>r�;<>������o^�;<|�	�.ۡǚݿ�������e`�Q�.:3��_T�C
̟?�_��100�_���ԣ� NBF&����V��H���l+�W���	��^��F���I�
ṕ4g���~j��W����I��S5TO��  �rV��`���:�D���EԀC�r���Cǀ �[J
��%p]ꌸ��賄\��7ɖ4��w @ �`s[M�)&M��ڏL��KJ#�!y].�E��G��q�`\��)%�z��& $���x�����<�-��ޛ���Mo_S~Qi�_�5�t�^����s���W�
�_�J��'Z��p>��ɎWK�����
d�wYTf55Q�ѵ�9mj�%�ZF<��������@S~�oP��̅9!����.���O`�+#�z]r�mV�$��c$�NL���M_���cL���~yr���p�����%������ ���f A7��*�Rϟs@y�̈��/��<{]WN�L�Z��C��4����~��h|�'�f����2���	(��|��8`uc#(V���ҿ���_��ל�i���ۃ'��y� Ѯt}�cy�� Z���3̕Ax������	5��2*�F�����$��t����,�8�?DެEXN�dj�$%�1�% ��I��3g7�:N#��k��S�^�(V�020�f��a�T���AA�+����I�YV��(/R`�����Ŀj���)V\I0�m7;��L;� �)�"����`ɿ����g
�߶FRh�$X�0��qb�V����F�oF3W=_?��*�.	�J!��Ӻ�߷I����T��gR���X�@;F'!��؀f��'����!�!#+K��p��AE��ŗ @̋^�ߞ`SE��i�e��^�ln���K��,r�!2C[�e��ޑ���9̟%:�����l�g �RJ;r,&QIIq���h��Q;2�S��/�.I�c2�N�H��T�_��
�Z��05��u��?e�h��� ��X���?]�γ	Vv�/<<��������#�w^�������5��=c��'�T��?.z��)�'�u�T�H淬O��)?�X�p���O��D�peYYk]�T�H��pKtj��"a���-F��h�����o�\���$E�����p��N't뾔�:u�����Ɇe����<Xu��ϣ���h�oDJR8Y��>��(�����m�KȜE����kӆ�����Gs�!!�)��}q�=����L2��9*�����h'�C��� �k�n���3(&�26��Mu:A,ǋ$K����˟�w�p|��O7E-C��x,7������d%B�W��+J��$2)'�%$�����:G���c����ש9Oŧ�		���""��8I��&|}	������:�:�D<&� ULV���]�ps��5xu{�65����R�����Ǐ7E|�ױ�<�}=?�n�c�.��?~+\`�aU��Wr�uY�8<N��iP�H��$H¬��;���&H�ʯJ�:���,���.ڐÅ�<�?�3���T�E��/T�BsV駓`�GD�1؊QB�C t8��T�<c`u�����鲦k�i����W_�gG�a���K*i<D,����`;���.�z^z�l�MWV��3pu|�t�����C�{�������n
��f��8f��H!�;̣ۙ_�M��:��}��J�����k��O'�rU����6z	K�^^��z¿'p�"��l,�^�R� �N�G~��E��s�fPVy9>�ŵ�iU�\�p-�;2������ں#�U���lr	EU��M~R&f�������-'�������V����ͮ"�|�����v�P����zLk����J�&�H{JM����2ޒb{��{��VY]�HHH���J88p���;,C۽�L'��H���Ņ�z`s"��c"3+��R#�l9�g���Or�󈊼p>\U�8m�{�~ _^,+�?�mʪ�P��,�[��X ��-���5���s���\�8��u�C~?��]���X�@�n�e���	��H����bM�����22��ǰ'\֮���KGG���L]��y�1#�e��t��VVҳ�}6�6��&���#�ͭn�=����L9=3�:���gZX�5088��v��I4�
����}7/�_}h/��-|K?ЋzzvK�hGG44Hr��1�5�T���>{4y�}o:)-����G�8��Z�
q}�#Ԑd�l����� \IGb�J���t�nGo���g@��1��V$�
�L�.��οy�<��r�����H���S*��x�����U���G��W��k��LN0���)M�`ac�R��4�F�]�ܚ�f��o�5��+���;>��X��_�`�_�%��x<犅�E�c�!$�%��>l#���G��|�V�F�߿ӓs^�W4^A�b��>"`��@W9��v�ω�Gz�\����5�qh�<a��k��.`�jC3�;~�[��Z�D�>���ĔOc/]�P������J��r��[Y+Ϲ�SZ��@2:/�>]0�OUJ6R����<���<)Z�{{UV-tw2�2I��okR?��ea\����%�^�!�����������i��h�&���`w�V����L�����v����3���&��o�]�4z����+����E��iƓ�rL���*�Y�a|a�~��c
��8�����uh\7�����9L]�@ʜQ�C�F�����n@�ӯne7S�Q�/j x;��LG v�MG�
[j7����K��S�i��]JE⟲d6�s8�e�Դ�3�a�	�#�0@	~��}�tqi)��t%���"cߟ.������N���o�ν�gmfƴ�&�ǧ���M�R��[8�c���Ңy��?)�v��@q�M�H����Y�ϴ�����<���H�u�_����z0��W��^�w)�RW�
�a`p��G<�(o�Ͱ:�d�����=�,��0 2�o9�����?� *�H�!	+<ȉ��N..�@4�L�k���t��n�������j��)*y�B���h�����f[d�(���ʽF�P��9��4�}_�\)�>sL�	���O�t�ds3�x�]`D�]6�[x��ߐ,���o_s���������77�r��忋�1����������)� 6�M���L=��m��s2{�A-й�`G V��.&&��0��L�v;̺:;9I<�*�JTT.#�<H�C9���g_)���h��Ա�{bVH�����`������7���iؤ�h��l�h�
��gH_��G�x�"�Z\��-��㡀o@{�S�O+>��#EB��J��$���%��ɯZş
�Xdru��a�y��R0)�G����LS�GQ����祝2��
 ۿ�Ț�o����U:-��"l�Z��K�Ԫ������ĂP�z{�&9���U� �g8��^�����n����3?���1%Ȏ�k���T���ò$���1�� 	��V���x3`A��ס�\�0nj���]_
�c�g�R>~�������"D����l�c�8�oZ���nJB����8���D�?�o��#7�#n]Pln�:��L���ޒ���+FX��L�#"�?��?Z��S>I>]>8�,څ�	L_�5���~�pņ(;�2�Vӣ&�@+*2J��:V�H/l�>�58��������7C5�|l���8��zc���D��qQ���|���/����E�����ɼ^�&<��0i�����e&"7�����{`�kHD�������aݫ^=��etF��5?x�d��vV���c��
A�0=�Fx��V~z�Q��*q����vo��hF}�+-�*M����ʖ9ϼ��}�x=U}�賈�N6-��//?��f*��k���f -C��795��&Q?���,��f�6�<X�n��.Q�3])Ȣ�3_E��/��x��/_�XVV̫w�%����I�s��K���&���LP)���N�x�y�,˹���Pn��Ryc�FTtN.1��{��qۀY��J-M��C���-��_X	=<=Mf�ҵ�Vb*�q:����[�/�n9?�d�}F���<NG�h��ae2>ckuub�6���)Q���?��5�Љ�S��^{���5[Ue�%�A��E4N&��n6�W�-К����;A��O�O� {X`�$H�D����q����T<���%��X���!�;>����rG�c�cs
~���/d�Z��<0��R��7����o'7�����ѱ���N�$�<���_2��#ظJ��z<����A�	@k�t��Z�b��ed}���S����ńVU^�R���Č���T�S���L]�CB$�yO�M�yz�6{�+�	!O�L�au�Uس&�m{�q�/k������LN7T��ӼCϼ�g�7��C�{|����$�E�&���/�6�xM���cx�+�D6�>隶uX:������#��<�;[\�隧�{B3��0����D�)��G�R��W��5�L�o��Ӿ�/���`Q�n� �/٠`a��q�m�@�|M`cz8�1n�b LJA!++���'E���jQx��N�����i�׊�?Eǁ�^�o��E�vqٝB�ɱ���T���MO�
���$�<�Q�����? o�� ��lc�h�1�GAC��M����F����@E�\+}��ܜ�A��k]�7������:R��9����Dk@��ɻ�]U'a����-��[C�*��ծ�����l#��|�V���9%���c��97����Zbu��z�z]:9��������bŽq|\���~R��u���#lr,�(��C@�4�Q��@� ìh�5�*�%}4՚��kuqÒ�o����v],,-_1��'�US�}�d���aF:Ǣ�=R���I����*u�qD�i�)����HT��~"#�Q+��� �WBvC,�D8����=v�'��?M��~(4��6+u�v�{L��F����l��C�[�E�}����4�-� ]J#%��CI+!J3tK�)� 3t9H7�w����{��g����}��{��9w,	z���������{Z�F�������\ hMM�g���8,��_�@NN>�<$|�[�p����Kr{�ތ��߿̴���y�ȷ����?>ʮ�A[��d|�s��]�& �u3��v`��߬!���WF��)���u&�?�BR�S��o��/F�X���ϗ~����A������ruq��,F>4DݏY#>�E�m����l0��N���C��ơ�<�&�s��
߁_��&y�P�o�J<���!���e���˛^��s4k�5$=�\2�>�ll�%^����8x�����@�+��孲2����}���Dd)$��	����E���������s������𛡹�.%���I�4��P��&��EߙJ���쪭u�lfw��߂�b�9N�]��[Uن��bxM=�ؕ�{@CI���?�2{ޝ�D�K���Ej�ő$ ��p|fK�<O��K_���8�>��)VgT<�ᴀ�Qd5�6�$4�l��b��D9 �1�ސW%�b@s�I�tnS(z�7T������LT�szҖ�*t�T@��vڌ�=ʣ�l���� [��~�����n �X%L�k�>��Ǌsq�H\�.�D8?Nūl�8R��8[�?���3��	��c->���5y��\9�7�ʙӭ��IW�u@�}ʺ.�� �iUU��e'��>���$����b8B��;���5$����_+��u��(��#�[?G���@���h�0&�m�E_t)n�廊I�D]w�4Geů���ƨo=<�B+�]�H#�1�D'ZmkCa���^8,��D�M,m@ɫ�{��:�k}.�}�?m��d�]�6�����|�հ��3<��dj�on��E�ft&R�.ܩ�w��:�Pm 5��Y�/�rC�l�j�	;[K��^<[�)O��_�)3̝����O�����;.9&�eL��dd^�s�9;�[�`�S����Vx-�@� �f��>��/+�\ϗ��������PL(u����Tp(	�P�D#*L~�G{<���շ��,�^��@�Ɔ��i��M��RE	��̛t��I� ��[���h8�Ԧ���ͥ�s����v�]����8ݶ5G�ϱ���<c���T����1�l&����Lo!ks�L��Ӽgu�ߨ&�RR��ɷ6����[���?��P7s�\��\���rgtz4�I��E(�&�����Í6�/��[W��}�X����z����-�?�"���̘�{���<h� �+�YЧ�)�����جM��_f�&�����"����su����(k7흁���5�i�Z�8]Í� �Z�`1\���fj1�n��D���}8����+�<���q����h��h}��9��oϹv�bkro	�Uw��n�\�,>�����U�#�Y;j�,��8�����kv٦���$����Y�����i�T�ǁ���9���^�������s��OO�ȁ!���[_��?�y���&|�f�u�m�4r��t?��?%�KiFi�)ji����}���a��C�9o����7�)�����t��i8���^�+����ogƌ�"+����m����6�-��W��8��!��H�[W���Ƅ��k����y0_�,��.����Υ�߂i�N�N��_�=I��N���g��x�kGFn.��G��=�������(���g��#�U��Ͽq��3s����Q0�Ԟ�~����.�}߼�$+eZ�򤢒 ��>���\���QW�(��5�����B�fO#�ѯ���&]ߊ5�9��Fi�P�E}<v"�z��3\����B�k���J3
�)S�����Z��E*,R���dȲ���v?I%��g��K�ou���X���VA+vӼT�L9���?�b���'!A�;_6�2Z�奏�>.sZ�L�;�3Q�T�^!eFf��h�"�i��^0����~N^���ԝO��B3ߵ���@��4"����]��.-�5}�6����>G̗6_����:�
ǳh����&eH�j�<���5�M�\N�����T�O�8.c��Ɔ�����I�&�)C �s(�L�󁝱�2��|���h�*�p?��4�%�o�<r�\�܈Q����%5��4�m�^���(�����Iq2�
�s�̴��###
yQf7Y�yh����0����!S$��fd���M�ƛ��v�3�@O������\,���P-��響M]!{�ſH�V�Q���E�3r���,�jlb���@>ʓ�`���65�������i����'�Cy��v�H�M���!����������WT�VF��-��y�}�=J��u��&W�6.!���%f�J���f�QPPP�ps�(K8���~>n;�&��Yf�"�m]�_���7A�=?�/�
K��Į�����	��%��	Pe�@�#iC	0�ڙe�����m���©i�8��f��͓J���}�_��Ԅ���!�qݖK�/ɥ�8�D�X�ȫk�'��m��S��u�^s�%��.���%�'�K�s�s���U��؞:⛲8B�@���������3��~���s����B;Z"q�X	�Ӷz��]�����諝���� � ��+H�br�^����Q4oO��":K�%�|�o��kY�c���]ݏIi�l���fl,�ߧ�E{2��ߟ�ٵC����U�I�"�o@&,�s%�LM��q⺦�b	�ͱ0]�ڪ{ ��W����׼�M�,�޹ JӉ�3��>>�꾛[Rߣ����D�����KG���Z��c��� h���ς*�k�07�w���,��G���!
!����=C}K9�0Ix���#sl2W�CT,7�07]o��x&��_e~7�#�#�Xqx��� �O�	퇼A�x��C	��*�ʢ����<���Y&YS?چ^L)�;{��?C�u��H �JM-���}�\�~�A�&���ˑ�k����񗍈��#��"�X\w�hJ:�/�}����꒞�/��(�H�C[������R�x�B}jH�� ��6ss��trrµe����/������7�m�l��x-.� _���BJa�In-�!+�33����|�N�4�}}}�������a�����~{���T*7�~�f;?�1U�Aݷ`�<�â\qo�q����;
����;v_MU�;wE(��@I�����>������Vݯ-�܄P�\P�}��S��uCc����������>�o2��0�.j�H��6N�iu�k��PMyy4^_<�N�rn9(2�z��:U�31yr��J��ح\��}��P�����=�΂p���Ĉ�~R/wC���]k�MLS��
0����ٺ�UB;0����X0V����� ��֫	��x�0�<{D�Q-�cu5�L��8�h�p%�È;���^s~II,UW2�L"PACGDD�\�3ti)Kau���S�A����e���@+�y&�,K�=��m�������_k������ƾ�X���-Qed���G���%ѩ��(,Y�<����{$U�q��:X���gj2#��j��.m>�!�un�z��ʊ��>�eq�xM����9�fc�n,�_��T�#�?!����X,Q��k��7�UF��˔�$��%����Q�Ғ�w|pljQ�"	���26��nK5�kT�g�p{�~��A0�I_TL�5��)0��`m�0�^*��K�h��9�f��
��M}0�6��(~���)�z�n��Bo�آP����:�H�3�WPP�h��?��aA����F'��-�������n@��ӗ�aI�Ӎ6�y4'Vz��P:Z��]
FN����&�� g?c��z<J*U53�D���$�Ǿi��F�]1����w��5�m�����>kDM<��Vvv����\����Hأ��uѕ�|J�J�|����[�S��'3 ���������un���Ŵ6���ݾyu5Q�><�(@�P|�W���S����� �z1HD�B�Rn������Iv_�M���`-��f��Z�7���a�>����Ҹ����^<� ��uYP���ۤ���M۳��X��S'ee=�gD�{�]�V��,�o��y���:=�5w$�v�j�`$0�y`u��4�\���ɋಁ��NI�3����dd�X%�Js%%�d��j�A�f'�J��<㽭�b�����r�&X�MO�z;��h08�bW���93�]V=����=|����-�ѩ��U����!��L��Ѱj�����Jn�h�j�
��S���5�Қֲ�2۝�O8� RME����u���DӜ�W��<yhQ
�߫����A�5������u���Eǿ)��^�:��1�;�h�%���8��;;6Y>�ӹ�J7�N蜍� ����"c������nH�B �zJ-�����ʙ�D��9�'��ƈe����nR�����~/?�H5�&W���1�((W$�2��pc����f���D���i����KZ�e\\\�P�����1��L}R�9���+�:C`�eT�� �-�E�b��>ꚓ�&�ZB	j^���%Xe�I>�d�ߘQP����>~xܦ�φTvIMDFe���r,{�p�>���
D(�p��o3Վ��ݏ���"���1u
N��椢��7*1�'�)SX�(��B�|���u���gM�� 	��ܗ����¢���J�ޤ��,"$��j�N�N!y��}"���Ç��&R�7M&]�&������-2��S��%]]�i��l|����&�o��iNz{�����������NII�_��k{~hc4o6]1�� �kw<��
vV�3�;����Ť�^����sfH �{IQ%e�js�z?�iw�hH�7���V��+R�\ A�>�����;Pia!5O0{v׺������SHH�Y�C����p���{��"��/�^��X����a� ��99��W\He��h��f}k;�_�|�pܣ2^6v��/.63:�����*7�򑱟l����� 0xND$�"�g�`7�d-33�X�."2� �8[�9�]�Ƭ�2q"��)=�P/i!6Oe�c�h��cB,44�����r[M�m��4x��eV9��0X/Ǫ��s7�n�Eז\��L�B�����3����jj���M;hf�JEO�gPppLll���̬��D*��_�ѕ'�9kNM�3�Y�(�/�A�� �jc�d��`�?kw���X�=A���Z����ن�lD��ۥ��f���m��[��Z?��(l�ث�R����ԔF6��d��JiZ�+c�t���9� ܞ��4���(��
�P�E'rq�3<Gv���\���Ż���կ3�!�㠉56�]����-�*��2� ��r�*��f]�H��,~z��sx�:"5��k��ōI-Q3]�#�g���r�ځ��TS� 
�>�����&�W�'"�5/���v�1�̮����q@��\��`��$�E��K��[�(JIJ��9����� �[r�!Hk�0kx���h�?c�p����+����'=j�0�ag]"Wߠ0��x?�����ۋi�ǀcf��a������,�:[jɈ�?� O�����)l�������!�IC}�eU�*	�-��1��Yd��V2v����r	!i����7�F����Y,������r��cm�1c>}J�5,����R���ӕ%�1����R5�ç����ݯ$/�h�yy�+�Fc��w ��O*�H�%���� �8=�DG�~�ݖzg���?1�.d�.!Ϣ},I	�(!�p�H��Dg�<���ӽe��=�o�k����
GTk��x��~<�}� ai�j�t�p�
�����.Nb�"�Ζ����Ӻ�<zM+**�eT�1�U~���?T[�a� ���� ggt�Qf���K@����mj�r�D��<-"#l�X(����x�����f���9��~J>8b&�?~�;I o G ���w97@���>�Np�+��&k�Iu��.��7�6v�O�����O�3�4��z� ��������^oO�IHt����)Ni	�d��b������)�R�>{=�%�{�ġi��n�/������$!�j.�lk�� +�ߟy0�O#@a�z� /���ms�՛Z(���#:�j(�V���l��AD���{��մ?�]�K�v�a��1~�!�q�іSWd���D��3����%(d%����^>��v�����J�c��x��tE�g<& v�4±䠵%���Z\J
��`Ҽj\�$i�!�-]�!�y|���� N��@xxxbRb���i���`�� �bҪ�����nhH�:T_@؟g�Q��?�\���~9��B�����;h~i��ͅz�QC�v���_�������i��h2����q�e�mr����euu���y�Y_�}ds���-j\ i��*�4Uk����6������nf�%��Ĭ��<w�Ҭ���J ����m�h�������,��{��պ�h�V�3jd�v�gR����Օ�̣$H��I�3�KSD}�~wS�EbF4��h�?_t\�� �磕p������kh�I_<3��za��uo�I�?ѧ�{��"�	IfN�)پ��MMM�N�:8�&K��AaSeFLzMa�b_������ª\�HA�{ey���������@f}�:�т����N�$++KZ��mG���)�����#�;�q��F{m�aY�:@��@�߾�g����aL麩�Б��4���x[��)��B�w1{��s��$�s�t��/z�A�E�oE���k��<f7Y�s۝H�`9��M�_ژ����Lh���P�Gޢ 2L��T�;R�b��1��k��?~\A��ze�^�Y��N���tK/��=�B�r��8d�

K�߭=8-z��#-K�?P�ڷ� ��cfV�9�1��"�G����f��[�z{�gVp�K`%�:`/����̳�H�� ����o]���6^�c,¿%�9"y��kaʖ{�G}�ۇG��C�]7WH�zg?�(8ӺaGmpd?���"�/���I��-�{s�H����j��^�!@����WTt}� ddm��UGl��)��"�����z4��|md��� ��LJ��b+KKÅ����m���u{ۖ����9> g��ق%�A�A���lv3oXH�}�y�M�S��_�#汧���l�J�#�:|kL�I�LG����5�a��\I�o5�C�
���d������]��ze�5�Ch�!jm�L�4�p��t��&����y�����w� ��Sb��"|�Q	]���'~�SH�*-e�"ڀ7e�f�zR8�ݑqsJ���Q��d���pG��X:-f�A�^!��A�-HM��GǤ�M��z��YL�&�
뵔�tʊ<�/�ِjC�A�S�a�����|�m��a���Z����\ua��C­�88IVv6�y�u5�ϹK�C���ЅU-�`�~��?�*7��2���7*v��fq�jt
bBo1�Nh��"9�MY�W���|��<N:�~p�{%A��ђ��* �^<1��L��x%F��)��K���a��,�`�Z��m��.�|�� Ӟ�9�|Q�$/	֜��n�I�ش���������Z�	���КpN5���*�A aʎt��SN˚c�o
q����g��S��U�v;�g�� �W�V�̷5?#��'DB"�WJJ�q�}τ.��ԝ���x�w�|pnS�������~gxV8&�5�O*��.
<�/�$K��6���� e�M��}�����?D��/
6����� 4]cZ+*.^��"&n?A�
�"���,k ���z�և��gԤA�C�ƃ9+9�*][߾~5�Y�$�;i�i>����@k����w��;n��D��Ԓa�t�
������,�E�l�vJ^.q�>ݫ `���qr�v5e�6���kĝ�8����ʘ �%������<:5�D2�D���4e��1|1 �(��w�YYt���_TJ^��VR.���+)�I�Ø��V���F�+=1�sUI��� Q�%���$]8����0gB�Ϛ�DIt��5�����B2	��PX��ݻ������lR2�A@�#.�|�0�ݜ^�{�ϣ����@��	�	
���|ך�%���� ���%,����A0��ۋIS����0V#8M�,�%W�߯h�ס[�柝٭�G�޼ys�ڽ3B�r�.G�ܐ0B��U�Te������Rd>�ŚS��K����G	���C>�@�$CR_cROY��5�I�n�+h{�)����;��3��6D��(Yy"[���1���5��a��)�3�����B�X+u$Rx�����# �^�sr�$k(r0X�f� Ar�Ŷ`/s2�#5`�,�n*�s���O}����md�5�#�|����&di{�f�m�{�v�w�_�6��/̈́p���v�.���7ɋ������I�NMEq�ջ����.|��;�:�'#7���Z��#��S<�ʮS&����73�0�G^V���N�P� �Ѓ�8�_QQQj�i-U�GO =����:xai��p��
|�H��T�0���)T�[z�N���I��ӫo�b���䑑���ҋuQ�R���TYEeT����:Z^���.��K8�]���WW;�GK;˜OfO��䩛&&���Q���n����}[�!  P�U��Q�_���uqqq��Ɖ�����-GԹ��"=�q��&�5Q�69\��	���OZI}�S�?�]/bih�ڽ�&̈́8��o�Fj��h� �R���э��6޼��B� b�e�d�|"�@����@aAo<��nI��W�>����`�M>��JŜ*�r���Y�lȢ�� �g��f��������Ȥ"Iv~t��6&���kO�L��o��?�v8;;���^6���6;#J�S�nS8��	jaT�
|�O�}���I����C6�0��S�o�!��-�Y�tp�z�M_Zf���T�;+ǚ
�c?�!�m"�IS$y
���i^�5���}z���-��ȸ��[[;, ��R\��QFAfX/��1����W,,���V�B.���*�<���@�z���׻W�B��PQ���QdF�����2�K�	g�>DU]�M�D����M��S�P�aƎ|�Y�G���]�.�K�� ៥���u/��e�q��?$��������܉ ���\����aZ&Љb&\��_�>�Χ������eނ����U��?���~S涣}����(##3l�p�G͜V������cW�A��0��P
4Y����k\9�K�܁���Pc���6���_D��r�,_4g���'ge���G���U�ǿ�?�?�n�$em�*��*bH��xX��,�ʽ���|�Β��ם�e�q��z�[GH�KU�Ϯ��i�,�d��=NN��:��K@�(������-� 1���阵z�)wu��
pL��d٥��A��.wޯ(�w�}\�����|=�yG��Ԧ�}P����m:É���g�pq��:�_V��WJ�fm/;;f>>"N�0{g�aT{X�9P���f/�1�����90�&cf5v�'
zp�{� k�I%����@.��&��j�D�S�K�:]c��㓞z/��ЍR���]Z���sk�c����R�h�� �Ƕ�	��.��km�1c!Tr�W�N�V]�A-����9] Rv���_n8 mӜ �l�� Rt�F'������bk��i�H�� �f�`6bح�x���+�)L�A��s� e�E|p� ��񔊼TVl�5��խ�"u�Nm��@�燨Ҳ��EE�TۄW�@I^�W��!�'�#-��� �u"����~T�A�_�+��L�W7,���B��@
<�?��T9��X{BJ9N�<��� mSH�t�p�J^T��$����K��PAA�&��}����u~I�����an�����5�P�}���P☋�5A��Ky�Z:�'r�f�B�>~w� �&��&Y�׾��s��h��sr�_]�p��M�/���np�~���f`*�x�<D��������bğ(D4�~��|w�`�F	y��O /a��	������-1�/
o�z6I ���OCwxC��<{��|�Q��݉���M-�<�`�wZ�UP��1���08k��J�|����Q{{###Lr�����8�t��!���2�+@j���\��D�7Y/ܥ��
��KH���_[)++?
97�튡�<'��4Bh9�2z�p��Lm�Ti1t�lJ0:�*�B�Mq�-�1���fXcJ]�6�b҈��2q@*���Xc>�2�O�6Xt�T/)�#W���cl�~+�q��V��'I�|���naT#�O��W8���<vW�q�"�j�����J�Y����;Ѭ�,�o��QdH1�>�F&��m2���GMM�v?�"��y�?�G���
��w����Z��?qtA�F(Mkk� gڳHG�*\499Y��%���*�s��v���Um/i����w�&�]�5S�����A��k�+���ԨMG^ͣ	���9/d<0݆� ��T�ed����I�ӯ���׵�������!��}��m.v���������n�U��ycm�₻��^�}lF�J��a�� �NWdLl�H���j)0Ď��Ё��%�U�S��3$@{@�\	em��� [�d]�����]r�ς��Ε�PS�n7��B"�t_�
X�M˓��V��#E��ݾZ���Z˺�_��ඖ���y?[����+N��a���90���;w+�z�"�9�.\�e-B����z��>��<��V�)��bzLj�̯�D�;�R���^0���zԻ��!�@�bg����3��zq9*+g��Dn���� ʉU�w����7�S�( ]�
Y�� ��qh�1�>�X����-{v">���<�?��:QVW���!�镃o�Ȣ�^ܺA�+3	�-���8D�m(]�_����?�ho ���GmAء��,�:YS�����{4�v����܇���R�lO��r�S�z+#�	��nGOI-������ǫ���~�o�Ó0����K�#M-�w���s��Ðξ���3�c|�z��Whooo��Q�R��;9���6��(���_1��.=���
����=��쥧G���A��Z������w�h�5Xb�������gR�~v���q���\c���\-��5��|�:�a:���}}�LLaF;+��T�#�>�>�Yk+��	p�-&���+��s455�u��^�6v��RxC1��h·�_�`4�=dџƃ���P^�ayIm~��������{��7,�X���p�3B~��{g.�;~0�;���b����>�:]�۶�:�/j:bVn��: |��������醤�"�E��Ǥ�H���)0���P'�׌��l��)�H�f�� ioK�:H6?op���W�\9
����çtDx/����y�'��z�xtmm��&�~U�<�~z��f�1P.�KZ�`��iJ�{��J�*y�v�@&b�}	��<��	Y�]� A9U�m����u>Gp� ��z|k��'(����T�.U����N����I���#�} �))[��(�>V��<�7=zJ�ܵ�F��4S3s�Z?�����=��U8�J���-���$���̌�)��J��2�-������2��H�m�p�j#��(��z�d4F���ͰN`�p���Q�W���1�ߙ��&U����rw���ٙ��f��cYST�\���Qה�
Y��W�gF���y�������VI}��O�3v�i�������/�|�� �I��QiI��՟�X;��$�\�9���!AH�0]�_t�{w�����t:%�LE۠�|� �)(P��L���F��0l�^�-%�8���J�m �������'�>Tl+���*k[�3��v�4����W
�Vw��	�a��߾�ƃ##|��e��u��mr �>���w�*;�'��6��>tvX�v� ���;PŖ� ����������� ����'+wrb9 �����0F�%Y۬o���ԁZ�5$����}�54���6�ܖq}ڥ�n,p	�ĳ���C(��&�����ڮ�m����hK9�|�uq����>���% T���U���|�k#!�B�mKĖ�����p6���sr�]����"!������jq"7CW��.�t�2R��d�]��?m~-��h1?�� �y������_�~Muf����l�������%�x����_�NNL�Ӓ:�RP$����{���������8�~E����"�y䞶�ړ'�c�Jp�f$�BC�������0ߞ���zx𡠠������ f� �8Z��
��²^�%��h��$\N���9��**b��d��a�K@ :��2���#�s��t[����YF�hXK�����9��P��`�5�>���|:���)I[ML�= �v��h�������~�@<0����h��� H��D�3���$
��٪9ښ�N��O[�i-gB G�CP���m����{�$�')wD��}F��j�j�<�^4"1늤��=��ha��w��͞W��.��ڛ6����Vg��[��PW���\ZZF�R�|{��ξ�:=R��e�О 	yt�f�(^��Y #&Ќ_�������7�,�����K�)��< %F?4�B�=U��Z�E����<���9���B����������a� vX~�Jx��'***+�?�|,�M��U� ��썄��F����K�eߔ������-@��!7��{�c��4�
��ߡ�֮�`d�M���o����!����67l33���N+�/�3=����{���U n�xI����g�%�4�;�ZR�Z�	��������qS��G�pwխ፹u_R���Hy�md�
ZY+K��/���o��h���陙��H�&�<�m���r�)�r�Rtq�k���8O!�`3��_16d��p���a�m��}�oFJ�"�������F&�I������������L1����<Gr"�����d�{�<ݚ�4{�z;���K���g�=}:���9r�f�b�R5��b0���~��`���]�TOO�z~z�|��v�c1�<������ifΔV���u���O}&��	��G�<�k�*'Y|V�k��*w���&]��TUx���Q&Z��Kvi�P��[ ��4y�]�o�
��?Y�bݻcwf��6y͒��[�w`o�L�3���R.�0_�#�׊7�I�D&1s��l&kr�.	�|�Hž9�N2��6��Q��9TRNSXXx{��)%��֠�N+�*s�9��O42��\1@c�S��R��������VBS4h�ipc�	�Ȝ5w������)5Mi=��������Ղ4n&Z��	M�I((�>MM�r�����U^;�;pȱ���eP�{NSr�|}(��K}����Xi��E㗦e����8�ց	����L/lܻ���\�����8�B�f�i�X��+����=�y����h��*�zu���S~A����n��ay{��v�s�3�����&[q��v9:,�.��P����M���L�q�������K̟?�K�'�	�Z���L�s�9p�� ��Ɠ��w���1UW$ivE��˫\�Z�um��Z�_iմm��<-�TC�m�N	���٠C2C)v�X$)Oėsϐ�����_����y���'q�pB�����x���G�o7�(
��N�]�=<�	��o��m�s|�A%W���Jԅ�x;�"�b�Rw���#W	?��^���'33����u	��/U�BkՌ7al�+yl1ٺ��>��
,".�����;��0�]����c���Zb���_�`�/_�bd�!��P[��2�2}��C�R� p���ڪ���L��*��!c���w۟��$���KB"��B��7d_?~�վ�DZ��	pY�������K�M$=T����!dYY�W';��́(%7 >x#ɐZ�Ѷ�C�tf;̦L�<������NGʻ��/�s,p���H*F��\��V�&	�c����3Kj�Lr �#4�m@�� �9�婓�/f���͕t~W�<�_��(\�¾�a�<�� �~�"����
�H����r���yV�|.�i ��=k�'Ӑa�&�和�I �zN�"��+��R�G��,v�Ywl����Ʌ�D<c8T/��;e@<|����ȳ�Rו<$��o~�狭���!M�,�&s�'���I�,;x��+N���S��3G.����� m!;�������Php�\�`�EBB����p���� �$60�Ft$�ӟ�U�Ľ�̓+�%I��i�^c�n2�������# ~��ܽ�w�;c�����=|1y�^���h:���h���&�-���q��M,�3����t���3r\z��K`�����y�C6Zw��W�+@���"��Zd�u�M��]�,�?����f/����FC���h�s�*.�T�c��Kx�ɦil[%���0!�Z2�k�
���{�D�E�P�H
���{�t�O]�������~2e}��\��^&�v\H[��ޒΨ�Y��A�E���M�.���;��KW�mc��LȦ��2=����3����u �00���"َ;h��d��1r���۞���2a��@?xwe�H~�4�?q��>����$h��:��������i)6��f�j�ouR�����.��/_n�W��(����$�|��T��+��g�O}%i|?���ԩ��xH%����}������w,�������߄��Ne}(~�d��VTYG������n�A~��n�����Wa�Cz�-svX�������GD!�x߬���]~�zR���s��8���o5׼}��W��׺�	L?�۔�%3��ŪOr`�9��mɬ�c�t^It|�BiS`��K�����JW��3_Ҽj}�.qT��QT�Rq��YO猡���첣Z9p!;ѷOP���Nr���5u6G��Ε�ᩡH��%h�~Κ���j��ӳ$i�\q�~6�@b�[��[@K�қ9DUK�E.e�8�v*O�^��M�L,IE�o���r������Z��?��4c����=
Шч������$�Y�SE�l_5e+�HfyJ}�:��z
�y��MB���l�،�
�����b��dT��Mu�՜�?�O���m��Xn[w8�[�����);����CB�z�MBz�Ǎ!�R��;o9_	8[��۲JY�HZ���
�r*��;�����H����W����=�H��wG�	bU����յl�o��^��X��Z��x� �3����=F�Ѹ��Ϡ�&�@3E��3�^�l�B̞�q���)Ҳ�Y���"�(r�Y�/_0t3b~��䛄��̜�� ��O������:
�rč)�c�~�~�yA�+0�c�-'��7(|.BU��gO ʣJ:��
�=�7�	��٩`-���%��aYA��?6R��x���V�����rz9�T�=;�Bv?�c���x��/YvHH����k�St.,���}B����a�G!J?UgYů3�_|?�Y�������S7���CA�o���-\g8�L��/�?	���΅��<�9���X�����=�t!�׭�b�"��hSNa�͞��ZJ�j����R^E�4������?�_��ؠ~�	ѭ%=��]a�3�ښuQ���f|=ğ��B����#��+Gr��oX������cBeТoZ����O���`[W�`�"�{QW�)��Y�0lAZ��!'j���r���� �$
f�c�Q]���a����|�N٦F@8`ў�$��1t�2�������},��x��&:9ԓ_.��2=7BgLz\k�F���B�ޱz�̙�QP}�}��W�wG���RE�_�aD�Mv:�zD,�v&y�x��p��YC�`��H�lԵ���g�kc�����e]�.A4-C����TAm��K�v��+a���Z҅�>�:t���;d_���8�3��\J��U2|���W���j�k6�>c{3��3�s���ߋ5_9g��t?��#f�\'�'aQ�>��X;T�%���-����_+��9�@��)h@�h����Ňs���:��_�>,�~*����ֱ�Mt�w��Tɼ���}aU�C�&�~�&�����C) z�{)�؂"覓_J��K?Y�<��n�+<�JV��nN-Ϝ#6t��"��O������~ې��k��p��5�I{܉u:���������_�I�~*a�٧a��E\lG��Ov��n�(׿��a�-���)�(�`��iqNg��7¡���}���x@t���˛`������It�"����C�=���i��g���-tey���!�.O#~�~��Civ����l�A���5lrԨN�0m��]2*�nv��]u�c�6,8��p W��?�
�NV4�K	��& ����@ڊ*�s3�bаN�wXy��۽RG�w�>��6%�!��@?=%�����6E$LJ��s7�ps��'�P3ܛ��#�'
H�������κ�̓�;x�8�G�����ߕ��ޕ-{��S�Rs<F�s\�}7`e}-����y�]�����9�e�2�ݼT���q��sx�ﮗ��pd�NV�J��Eo�{�&xo���ܧ�Yp���]&C��:�u,��~�y���$N�?`���뷀c�\�n�}َ`Q����Eb�z]��_�D,ظ�R���>\.+].G���.���c͙r�P����g�ν2�uҟM��n��<l
2�= �
-W�V�LN�s&u�x���9a�`�Y�'���[V�i�Cv5���r�w��t*��ldMFE9<�Z�+��)ص$y�+��5��p�P*��D��D>��,�屋s�u_�I:tk^�G��2�
�t�'-�#�(3�}<�{�_p���N�a^d#ᣗL㜏�Qv����Gt�
$j2)H��F�y�Ȯ�Gmոx��RN�5��4]TT�Ӧ�[��[��E��nX@B���s��k��NAr���k������s���}ߙg��y��g}�$��	�w<;�z��l�j̆���[x&�P���q�"h�Q�lV�-���i��zD�� �8�TD�~>3-J�N$���=���ر1)���A�$�SX ��˿�$���-6���@���e`Չ�l�_GI�L
p�)�+y���-C�
3Ņ<��.�����m���Jmp/-8K��m��~ȧ��aL�X����sH�؋�m���P�
��p�oLw&[�2�`��);'儓H}OB[
�ے�/G+��&tXc����d���ݹ�Bf٨|�C&M-;��ь4V׾�A��%Z[_��A�B�0��r�gf��b��݁�u��c��[޴�@�%ɡO���E>
��ʝ��j��I��PTC�>�oAR�		��ێ�����[È����(|��Zq|��Mz�~��?�՞�fм�U��"c���۟��)N(��_,h��cP��r�?�d�m���PӅ����q����=�a�^;��P#�̚7[YֵھW�`�8�]�h֊��p��վė���j�9%���N�|sZ2,���@�'��\�������n�����<��Q�+�D��;�7��$}�a;B�)�:ԡ�1��ykn?_N�A5���x��利gE)�>h��D2�P6;4�\�(�f6�����S�^r5!>-	 ������;�����P�'lb)�w`�������oú9��4��I,Do���K�D���t����ۂ�s�9�O<؂��+�\g��xl�Ɣ���#�Ka�-�^��Q^8/{��X�!;y�}�H��蹵��702"��]��^6�1ّ)Ϸ�h��1H�0�P��-�9n���PY��O�B�؆��U��|؏{-8�K�S�IYe��#���=5m�C�r�/��k~�Z�+Yi̦`����q��b�K6�ŏ�JnR�y�<�e����;�Z���R�T�*~�btn�:P��B�ō��`'CU�fJUu�Q��Y`y���0�H <B�-$C{9d��*���9�:����zU�(�_��j1�'O�0�����ե�+FOB2�b����o*����&Q����n��sL��c����7��C���8Em@ꦫ���#��H��.yd�%Cj%�R$��F����J�qg�%! �j��-��7�	=����(OC/_���b�`Q���W���߮$3�A�1P0+ի|�S�FW�L�xx��*�|$�"Z�,ZhC���	��C�%���y}�d'����-W������`-���R�6-Q��
9�{�:��	9����/������U�W}
��A{�H�5�]����#�|Y�%K[���(ӂ;����2)�|����2��$��Z�U [�_�" 匟<�v3�������^!�	t�Gx��8<L�D�}6��'�n�GC��������C|�0��|!��n'>��,ݵ�7��ѨY#������[j _��H�p�����Ve>�������0}�2A�({�_n]�(|��l�W���Nq�Z����t�7򃏧�æ���[�#��<{�I�t���S���J�z��_d�0��o�f����e��,�}?�+b�%&z����O�Qr�$��j��^�m�-)a:5�֩�%ke�G3:m��^���&GLsA	��0��~�rg3#}du】䴧����L�i���̘��Z���+��Y_vJKҏ�n���BD�Y0B���>��;��<���0'��AL���`�jN(��V������jO�?x
,�]0���������7��(��9U�i����'�s5?|fС*��Þ�������9.�5�=���^ujF��.�ӏd<l� �u2����'cIai����K	�˦�N�F��w"�����L�ʃ`��`����D�e�~ZC��W�`�IE��f������Z֫�~�7RG�R�)�L'n���f'�&h���s�%灑�u��x�Z�*웭+D�i�ƓP���\t���u5s5H�M��O���ػ_&�NW�5����O{��A��8?��K�s��ܲ8�"�!PT]��A_s?*��3u������P����ͯء��Q-a�����& /Џ:���s�ܮp��<���^������	^���"������,��c��s��vۤ���|�o^�E8�m�@b�|���j��>��8P�)b���ڨ�uk��1g:��nJ�-�L.�����m4@X]t�t����[Q���:���� P��~*Ȳ���O�o;�W�K]�V\ۮE7��n���( ���Q�:��S�k�ж���X�ʠھ��/�����(U�Gu�-�Z|�ߗF^X�'-f/g�������O.O|�,� x�����˲����tx�߰)���L_��Ը�<wG<�"p?}Q#@�C�l|�%hzg�Ӥ�v�7�����N����C���Mg69O�V7�o�����ȳ��4��8���k��hG��6�&�LH��D Su����=�F7���r���M*M���68v�TX��R��H�xZ�P����Qp�.�LG��1��� ��p�ì�?X��@�`�6Q�0Q�8Ii5���ȋ����-�En؎7&<_�`��u����1��Ca�Bm�h���[׹g���Q������Q��(_�o6 �mP�\bP1;eN~�c�#���d�w�s��_fV�J�6����[�ᦽֺm�*r03tϮ"j]��v�)�3jM��w��;�����)������P�*dؙd��-��  ��޸�7��\[9e�Z����;��%�d��I��ΕN��!�
�+P}��ƿ�s��ac��?�i���9���u��%w��C:�$�H��K��WK��	T�B:�bG�y�S��9��C_������~�*�{��=N���\�,T_��4��bG��)<��y�	�ge�'d�sf�gi��1���κvp'�WG:�(^Q��nۥ���8u���#ԁ�O� �R��;0&�X��2�!itüx@{�ite3�l�#%s����Ȱ��Q5��K.�94���h"vq��!scۆ�?�����(�����p2��D��i�"B�8�X�M���ػ�k����(�����\�G��L5�A����r,ύHD���T�{�MצB0��Ӯ{�����Jg�����zя���%$���L6;��p"�ruhx�x=�z4@�Jn�e�g�E�`m��_�o��b��L����9�?���C?-�Q�L�J�r����8��hŎ3}��"�dNi#�B�|��Ť.���l����`p�|�������Xg��n�#�|9�����2֢&��c�1��Z�,�?�Q(��-��ٳ����ܱt��ׯdN�q��[����K��������x����m��o��DH��)К��q�}{�\~�}�O5)T%v���烋,i�*qb{ͦ��VOD\Ju��k4B��=m�
�$��oj��*��<�k"x�M9���~@�<o�\>c�,��X���͠�E�/���Ƚ�ݘ�Psם�����g���C�xG��fsh��
ѥ��ޓ����D��i��H��"�G0~����IOL�������T�j22I��T��j?c�����$��p�H��r�A.�D�r(c�
��ӯ��b#I��=3Sx�vH��jB���*6��y� Nt6���UeI��[/�G=i{���bzumG(����t-�,a���gAhll��j� :US���K eR	LϞ�}��N���R���m��W���K�\�w���J6\�O-��ld�%:���N ���dIKm��^ r a���x�,Hy]�<��=W���Te�>-N<9C�&tv�*$��N#\�,`^\ZU�&D����� �>��H&C#_kGњ/�ueӥ�XyRE_�M�� ��Zǣ��j�S���>{8�+GU07���w�1��it��Te�����<�U�vF6���QxO�@�!5�M�[9F)�W_������mg1l�� ��2�7�X�z�n;��@t�le-�=8�baa!ۼ��:�?2IOI��=�\	S�ũ[KhE�:z��٘���2���R�nOo/JL_��~+���W�(A�/pw��W����8vQb�����S��w�] O>>��:���������`/,,X/��������x�KU�%j���mK��D���q۟��.h[89��^����ë�Vւ�НW�G��}ۏ-]]����c3�	�<�_�/-e� ]�>�7m�gK���&@����������h>3�%�|S�(Y�����S/��ΣwN}�����1�ww?����(�]�p\�`���-��8R{��`F�Q�G �����v�{�(�R����m�����x���'����r����J ���/��+B��gmW�B�o+�;��-\N�|�K{)�E�)��8�b��j &# }��jj����7T��fwӗn'��T!� ���;��n��r\�/���wq��m��^�ڙ	��Y���`b�N:o^��t�#��}��7� #+���⢠�}ݛ����OT�����v�\exV��$��|#��G.�1T?��V����B���r<'
Y���fiBo9Y���-99�s� �=8Y��y	�l����y#��t
�������苭�
��7��=ϧ��l�2F�/��U�!ɟ����{إ����� S�h��5H�E� ��g�(��b�W�9p*���+��$C��ͦ��?E]�_�)���K����>�c���{�.�ʳn�N�g�	*n�oLy�7�2��ddd�TƧ��ӣ�u��&@�I=�L��>���o
<sc��d��K���
������x�<��S�&�m���<��~1a�����f��CMʟ`�!�\��mh��	��� @-z޼'j����rӚ����3Q�m�=):��Iݛ7*ߣ}WCHם�H:�䤍��]^��O�N�~6��U�Zw���~K���X2W.�H��3��4#.�����ľ���`tÁ�x�tS�VFr������S�ɤB;!��D�D.s*0���e��y_J_O��z��c��F ������7]X�ptl�9�U5��. z�����b���-+��1�J���B�37I>�<����_��g����M�ŭ�7�sBQ�s�W�V�bg^�0�'Hk��7�l����͊N�UWp�߷�����p\�XdW.��M4��*�dN_��������w+2&4�5�X�+.v��n���^���XR����^q�D�0z���S�	��]�jo�7�2������/��ۧ`eJFf&�G+�����fw�}\�Ͳq���hoϑ�ٮ���*8��`�?��]]�8F͝ӣd>R���d��&z�&��&#x�a;q���xl|<�k��t@�E��k�튾I�^�oC�H�O����Z}��V��=SH�U��gzn�Xn�*�H���J������i0��?������9CB��<ʌ�2��'���]Ǧ�q9*a�O|'YG8Q���4$|���<�n��t�&R�fltt�� �Ǻ���?����$�k�F;Dk�w%�K��xuro��<+l��B��}/�fc�*�^�7XI���4*q��|`U+i�	T[v-x�O��h�4HU��&(.N�<]���4=� 3q�6L���q4����W���B�dz=��.*�:�<�Q������V=�T9�aX�kS��Da�g��h$����־݂2n���]�W�wzMC��Ԁ�XԪW�#��_6���?n5��,�5Q'���z���d(���m8�bW��l��OUk����"��:����]������Zx��|:�F�׵ϸ$]^��V�Ҭ�]���?�O�bn?�WDVN'}��Q���p/^
81��qj�j��>�B�rdzX͝���0m�?)�gǒ��3� �W�F��/�&I����%�E��h��p��ld8�����\l�6�����*#����L�4��	?#;{�l��j���;x�L��Z�u�/��^��gix^z�!����EEK S�������1n�U��7B�_����0ږm7���R|T��7a��z@x����%Z��(,B*���9W�.�d��/�+�m麑���Ҩ�YF��s��D)�D/��	̄z��͙ �%oD�~�~�B��aa��RR���Lĳ���* �>�̊�j �0�w����!�����;�&�)�t�����¨MO��m��r�-}�|�EhZ�C]��T����t��n�}�����~�j
�Q�@JZ�rr���������i�)>��	�� ��C���뻻�ȧ#ʢE��k�ޟ�̨s���rݴU�������+|X<`�2���W��F���Ȼ̘���5�k�o��O)S�����8�����+����R����L(�'�8\�\�sC��A��D�Tȶ7��-���UR��k�/��qE6,�[�����;���td��К�M�w��a�N�q`��=!%4dF��'��I�\��D��k�KC��pAm�	�N0�
���r���IQ�ׅ�Z��lR���7/�=i�%S���Vʎ�K�yz
L��c�٤m���
V���oE�ל��N�4��x��L$X�������dB�l�8a�k�0�:b����i`����VaI<"��d�1��!�3��Ƌ0��`/Za¤r	|WZ7z��AP� ��k���q���������'i�Y�B%dv-�^����5?�ͺv{w2A�m�����gM#�V�]Z�!�Z����@����$�����)ôP5o����N���X&���'��L{jI������8���`:C�
\�Bx �]f_W�U�C�q�P�EIҥ[S��>���+x���>؆��^��D�%3��T6�������"�LB;xpP����6*��PA��;��ቦ�2�y�|^�o����F�:ڞ�X/�<��Ѣ�!N��$�InE�p-=�	�}��6�+��f�d�;WV[�C��֛%^m��[���}B���y�n=�؃@�}ûR�?B\5����ִ��s������J�eM�A�ދ�= ��Ή����������q*�MG�vQ��W٣��e�`3,~�l�S�џC��%���_l%6nExb�����v*_ٮO���/�7�R11�q>}y� �(�0�.�����Z��(���_m�+�G6���H�/HUYL��iAXrЖ"�Yg�F���E�����&��7�v��B
:����r��R��V$��y�r0��Ɨ�}����E�
��a\�L��^��:��_P��X��˯��}��[Y2�W*L�.��F���<��VS[�T)�~� �/�f�� r��Ɲ�T��te��׵�)�(̘�+�䐡�O�8	����)L����Cz�`,P����)�F�/��7�������3s��,�����&g�� �V47�Ma1�E�i�B���m{{Ԡ�MB�^�:��4���]�Jrc��{یZ|C˴}"@��'��%���EX�~m�PaduNo�DL����3U�j�����!3
���7A��ږ�%�L	�Zo��i����ƕ3�I�i�o�~�����XĎ��^Ǩ¤�P;��A�i����A!CD����D�6��`�� ��&*BB���IP�F�_�eR�n��9�[�\2w����������.��,����MFͯ��^O�j�=�ɅL�M�4zEH�|����!ʪN&-
sK�*ˍ����k2�{7��h�<5I�cʛ�")��d��x��%�0�U�Wb�w�u��A���a��_�:T -ӯ�#�����#�c��G���@�B1�mY���1&�E��Z�z����2'�U� h���̯&2��B+UrA�*�����Ҟ�b����XRB	��'x��k�%���9�+��*�f���F�����;ftKR�7�b���'�DVɖ﬉�^'@���e[����hװK�wQ����W[2Ex�~<a�ƣ��>��̭UCdm�������]��G�.y����Ƽ-�����թ���Y���N���y��t`��`*a�0�c��
<Y+��6ֺ$F����߿l������a��=���Y��q�p�q�+-�r7�|�`�Ӽm��Y���7�=<^=��A�&����#>R�B�"7���"U�/�0�$�G�)5��hYK��@!Fڒ����ѕ�x���﨟��*uN���L���㽼��OO-j�|����Ќ�%(�� ƚ �ȬD� �>P?}NܰӓM�$ ��%���E�����E�+�ޗ���C��0��!] ����.�(d��hXNmv�F�\qc�3��h-�ַ[
b�Wx�:������O7�V�,�,5o��>����/���$�=?�����K�j��)��}��:�4�fqd�p~,͹KV�sbf�zG����)�Y������?�`��� ��PM?r-VR�z�%��/5��B��Vn�H��e�^Q��?�^ �Y�����;ȧM���I{c;�k=
�ڤ�U]��0t>�a���B��on��N�7��͇��F�~C }j7!@ �*k�B�V4&zT���oE����?�Z@%���̮<����?Z.�� ur�i~�q�i�d�љ!N7��^�RQF��>6��%�i�cN-w���d� ������ϭh�#�Ro��=�͘��^-7��]���Ҥ���E��ZJe*ޒ<�k]��9iu�z�8�޿VdD\��ή��U���aWZ���C��A�;�,��_�-20�A� ˘��	�>9󣠕��I�%L�c-���6쌸~���d�l��jL4`'�{��w�QL~�,)$�?OC��͵p�X�����d8S�D���03l�K�v�U^�|J�>E�&(�h�W�3>�r轓ϫ�B�q�J&o�Y6��`�%H�]����~!�����"�?
��ަNnu&����n��כ��p�b����y����_�*�ء�;� iQ����2)8l�lvĖ��#\	��(Bq���!�'V�%$�kЭ�����'��J����0�X�V���k,5UQ&���6�g�`H>�/����X�YԸ85,�}>*qCkm��`�?������/�bv[J�2�~�y�ٽ��I��_d�y0g݌�ݻ��Qz@H?����7�����ډ�����{&Z��Sǭ�#i�Gcfȶm��{B��_c�<z9��n>�,��e^ʹRL�ڛ����h}�0��JQw9#��~Id���kM��O��j��i�N��<�"�Г�oz�o�J�t}�ԜH����v��韩��h�*�M���RΡ�Zg%����p5�T;V96�1g����lVe��!���t�l�%|�1*<�2�����Cc��Q�!�Ez`R�:#PG&1�� ���'UdI�3�m ѕm���ӢD�M��2��QobG���&��������D^Q�5��~�P]Q�XS�i��q�;��[�y>� �_ ktV>���M�
n�*��UP����Y��ڵQ�H�$͵D9Ʈ������.C!XS��s���VQ681������}��o��o��-���;P��T���N�z)�5��[�	�h�O#U�Wo|�kl�Q�7J���#|Y��l�EIOB��1�oi"�g�� ȹ/��p��z��a��^R��>���I/��K�]�z���?J��$a�6�U�s>�Ȍ��j.δx�hP�m�Egk�ග`��5���0�ܤ�p͞�6�n�wO�/�Uxm�Q3ZZvk߆{���n6"���f�>sS�U1z�2ӢtYɼ���^:�2H�s��Zư?9�aWg,���D&P���H�8�pt����(��c�(�}�'�|��H�
a��c�(������n�a�����@�B�i���/��q�v�%#4 ]T7��[��i�r"u尴�B;/f�`��9�O-F�{�Ql��lt<R�2��=�H�4�	v���IT
��&�Y���OU1hTύ���춻2\UM|È���~�7ۧ�K��������Z&yI�#�`B=-A��Ĝb�u���CG�F�1�̘Y�dq���gn�#1�> �9o�}����l����&f� �K�cE�D=,���1> W�5;~Yy�L�k�k��J0��������/FlET��
[�cMF��ҍ5�
c`U��m�xb�W���x8��j�b��%܈=��H�$�%�|�ܭ9�~���l����8I�K"#�m��|�s&�;�k�k�x
������^�ۯ�%��1B��u۫v���$�_EӻE�)]�cx(���w�E���,S���o����-�JD͞��9|��tn�-�+�\�b���o9�Pe!�Xm�ޕT	,�%��6����Y��9�8����B*��u��UW4 ��s�{D4x�����v�ڞ�\���AM�8�/�-��^�M7]�*��(a$X�v�!��
P�b��O#H��1��M����șS�&?6lp�̝�g��9���?�n#ײ�{�{���͎E�A)BK�c+� ����%G���d����G�zz�}=�Wf[��i)b�� ���A�4�_!�� ����dΉ������]*�lU�
B�:�$����?I0fx�6<Y����n��L�w�l�:*|��0u�{=w�����<6i,T��`�F��b����d[�Ҁe=8���mRYY9��(���+�/L��Ok��m/�mE�Ǭ�Й��9oȊ�b���Y�W���-��]Ss�P��M^�V��4��^�M�k�3i,X���:f��w�����'M��<��Ļe���l��i6��G���B�(�E���5|�����M,]#�����/����E�e�_��43���Y@{�t�L�����u��
b�+r��Hp���&�bm��E����.�,��áj��C?^P��u��3Hb��-���[��������"���џv�\s$�(O'y|��>��=N���Ekr�p����ɼlr�{�l�0��<�����L�	?����Pk���l+Z�&��H>Q+r]c�n����j�22�y��ݗj��b�tl�iNMqy��Y�X	eǁ���qh�ם�OF��oҚ�+`�j�@*���1թ��)�b����qRT�������.mg�G�8٪,ߥ���3�_QG�uq�#���p���⨂�e{	}C!���u�ȉ���m �xbJ�i�a[��);��h�a۵i��m�c7�K���"fTV�N'`8����Wr��"�I�����9���������U�> �P��
@��s�¬��n���]�&ڮi��YzN��P^1�ɸvX��Ȏٍ��LK$v���g��m�k��Co�Nc@
�b��>�_�;:r�]H)mi��}G�$׋ͻ���&h��L&'so���6`I�<������C%�o�R��L�1��4�=�g� 
˝�]����̲�w��'��oI̿����13Y���.�i�܌p��0������N��t}J�lȐբ�;H����(�Ȑ�7�*����Iw7����&z�����jJVe�v)��� ��w�	fAO4[/%=wD�\V�Ҷ`��)�����~��$�C@��a�Μ���4d�q	�c�c!FЭ���Q���_fe�_L�]&��HM��������q�����6������|�a�����+pbӉ=&�:.����j�DHLw�/0E��	����X�3͘�VH�_�ǅv���3�,�\}���~Pg4)_W&6j�0�_��qd��Xr�����L���#��-�F���WD_��u<��h�3�Iq"`\��C?�k=�e��%��I�/��7����&�3n���ND��cKH�+�n����иl%�>�di������ޒ�c���饥
2�(���	�O���%��Y��\��B��6�Ԭ�J�3�?���,�ޅ~&�t�g@�h'!���ˣ��������kQ[�����R��u$��Ie2JYM�v����" ��(=����j��?4�lA�|�!��k�4��:{�D���������N���"�#f/���e�����t�~G�C��I�j�aKcgq��{���'O�>Hs0�ӿs�Sf�j`8an��U[�r�f�1�a~��Y_��a�u��y��#n%D�=E0U�>�2N��)������Kͬ%嶩i�S��e=R�.c=�ﳃ��!7�G=��uP�|w$�q1�L���B��(t�^񼔔��M�X`�R�I�����Rx��[z�̥�!������f��]l)M��J�������j!L�.]Ꭓzqc����?�k+��m��^��As�YNK�2���%Q4�}��{XiOmWu�x��'�qC-"'d�Ax�<����2�����Y�Ʒ�*�5���ɕ���Jay`�_��R� �0m�陙�f����%�ڷ��`\��Q1)���+X�������a��0��j��b�x�]�G�T�dU���^Y��C���!��@�g3c��s8�6�uo榺�u�$qաE)&��N������o�������Tq�\9<6;���}�c 'U5�#�M``�����l��l/>�
�	�����5צ��L߳� i����<�P���輦�O�$��D�CǑb����43d��g���vķ��ʡ��֯?}w���km�x/$�� �ʏWC'~y��?XS�?^7z�~>9��Ox�iW^�H�/j@�,llԫ��6O���٩��W|��T�P��5���ð/�j��� ���FR�*}E��8�Zi����N��8�;>�% q�W#J:�g4��.̏o(��+B�e����\|'��������r������T�^O�֛�5�h�������H�*�4-����IB�6^-�������f�u��zt]X�aH����;+&�=�6!0.�g �'C��u��"H��"�V{ǳ�g-����Ӌ(�n��Eh\p0b��h�M�6�J2�Ѵz�iطɈ��i�4v���؛Y��&��j�㢀}r���!�[�f��d�i�NY��u�%i`�e�JU޵t������F2a� �Uۮz"�,#�-�{`�q��PrgLk�ɓa�Nۀ�V��>����s����ݘ�8�Q^!c|,�n��Ϟ�����~[OrT�vȗK�,
�f�f�"�]]�`�J��0��w�(n3jt�--I����M��uͭ��,l�Wfx���\#�|||Y�pj�_�_�͒�+��WC�	�]�:AQ����R3u�E2�s�O�M��e.4o�2!-Ɔ7�������
��]��֛ogʂ5Q�$�6�L�>�`L�voљ���V<MAMm��za��FJ���"
�90=���4�^#E����*�d:6me�/�0|�}����<3�읜��i~r�������<�.�d���G"wƘ��<R�OT��v}g�W;۲�Ϸ,��� gy"��ZZ(�8MF�"�Ap�V������h��%���k)vz�Vs��d�#@��쪱悁�_�S����ԍ\����������<V3E�:�ǳr��r��w2�al����"z��]���O�x�~	P^���oL��������VQ���t��vfR���nD��4�af��G��>�p�J~��M�ϳ�}�CVD��ȋ�jL�O	�Ґ(<_x6 ]S�C�����d���l�f�%(�F���=�K��Vw��5(�� ��H[��|�yI������c Zwʱ���*5���^kw�q�����e�$� {�X�P��Cd������m\|'�=ҽ����f%�������[O�Q�s��8�X��'-������Jgk�u�,�J��,0��,gL��R���������=�&�m�`�s�u�\�r�:���߁���`��^��9����x�oP���H�fT���D���}é7Y��ρH8.�f���X�|�w���A�,��=7]c�?��OTe��J�[�4�� k�C*�Vh�y��c��g��)2ν���1;��9���ά�r�hM�Igo<믧wg+#��:����2LmAi%]��|����,�2X���?bۅ�?���+O��r?S���>�y��Sk�/^�{ڐ�{�o�&�X�>>>i)���%%%��g��;�ai�n�x�O���2޼G@1dL�[��^qHe�mP\;xD*�t��\����6XS���9<��a��Y練�l�` �[�����H|j��/�*��E�� �]8��B���c��yqi���[�/D����P�Q`��WG�m�&#�e�� �=W�p�t	gFڛ�׫��rY�3'&���V�9P6���;�6n�e�Rcd:��������ȯ�Q���I+�,s���I�J��$��P�ҙ݁1 0�I�90&��֥	j�?_D��&�F ��*=�� %�8T��t$W����J�{ӗ"쏚.3��u?�&Bh������3�������S���ot�innN#�/�޽������
g�j2���N���(N?3f725]�ja�e��i�9��^�|2u��'L�?�GÜ4����ndl��~p �q���I'�oQ7�#���2��!f��h��8 ���+'��r�Gx��R��w�2�ne->��cnZ�#\�u�Z�BW�jn�^*����<0F�����d��L��OG���ռ��>R����ٹ`�X�I�w���v|�M��1'6K��q�o�O4��hv|C�w	zw�	:���oXx~����!$�R���m�L0��&
�M�u�E�h'$���e|�`p����s����!��,��}��?e�\�8��9�Gkܶ,���%L�T
A�����͉����V"J�D��r�g�@�$)����Q�����7"�暍Z	Z	�H���{,;�>�פ�Y�U��p4T���$MP<��EZi�#��#9�-��||��#�<�^z���P���Kp�g �����f���Ϗ!������^y��秜����D��RY��!�͑3(,l�B0(Q���>���-
ɶԞ�w񛳔�z�zQ��������0�i�cZ�  ֹ�<��=�[k;nB1��Iy+]�z��Z�Q+Xks	V��-ϥ`Lį-vԶe��' ��.����8|�ԉǍ���7��>I��|�hfp7Q�:��gR����������ᴙ�6��ZЙ��O�y~:c�~S	�uu���0�p{��(؋��t�4m����#�٘�A�U<ͬ�KR��,�����]�#G���Q ��`���LJj;C$i�O-�$}B��㰶s$�����ťq���#������z�
�'�6,����f�x�kQ@GV��"�@-�� N���׹��Pu ,�ϓd<>�kɋ�l3���N���nĘ$�:?���p��>D�&>;� �E������F+.]P�}=���A*���N��iܖ�������/-`�T&u-og��+S=bPS�d�h�8�.���;�'���n>�>���|��<�I���UK�M�	��I�R�ژ�X���0�wՍ���v�%��4$��Fԓ;b���a��4X�64([��^P�N�#��T�)k�����y򽡦m�O"�8A�r�� }���<����Dĥ� P�/�#L0qho��B��rR�`Xϯ�}�����N���D�����nXA|�s�y�?y#���c/M�����fNO.��y=�ۦ��2����N����4�hD����\����I�`@Z]����6��fݱ���϶�ֆ��I`���BMH�E�0�,�^q��� �a1m
\�ȋf��lb0ye$���\��]�`9Ј�cW����iA��l�`��Da�e@� 1n��7�Gԝw�\A��\�@����`���"���#ğ�����s�8~���S�Wd�`���m�е�5�VVl��=0����=�a����6Ogiq�=�Yuu���s�h�Wl9(��2˛i��)@��^��9k��9h�1IL���6��(��z�}�0x��Qmr냭���bg�4�k䚱�P���Sd��{�q�-W`�%��f������z�sp���s����'�b&�jOc���uK:��?|�c8@Mj]o���=Z�z`nh�Uޯ�5��X��������^6��od�=�\�1�*mc�{����
�R*�����ͤX�W�R�
�;���A�	���ڱ��'<f��1\���_"x�]x�k+���U��YB �U�D⯶�Bqʦ�E�C��Њ:����7>՟��f��5�A�x���N�.���P���K/���'*�ZD`��>7�*����)�]^{� t(��P �N��`\��I���zaaA^t~x����W㽼���Q�OОЪ}{�+/���f�=%FY�v�t ^0x!;��ɕ5�G�:ŭ��Y�H���
o��%�Z�o+�.ܟJ\��dtf�aK���?D����*xǛ�Sˣ�0�#�%41W� ��zöS�������|ɬԣ�W���t��e�X��CW��k
U�y{��d7�<w#�Um�o�l�({v���Ū����х4ls��F_�
�1����$t�������<���������x�F���G�[�E���t�t��tww
(�� ����%%-�ݠ�twKw�߃�s�y?��e~��}�ֵ�u�Q��nr���7� ky?��\��%����y �ҝ�3�'�׳{�n�l��"�K�5��>���Hl@�8\8�dpݠ�a!�i��@��³��s��Z��|�]#��Y��	�;��vt����\m��{)M`=r�ѦKMS�}��,��5LVOVQ
!i��\n�-���i.th�F��T�x�G<K��+Wړ��v7�b�'MSk�� z;f�aӟ������n>Z��8+�8��{|t�@i��d��v|��I/���y��� �;�f�<��e ~ ��;��]�@H �����z� 鰻����&��$��1|��+R1D�6Ȉ�ʳ��5ނA��6��s8Mu���d��=3:�ϗ����2��E,��5ɺzZ/êl��'z���U�X�S�x���!�R�������_�����ta;o9��uH��vc���gG��1t�j~�m C�
[p��Qff�M����D�0�	5"�ᙡ���Q���H�	�A��Ѯ�vB��������F�Μ9dL<a��*!*rǟ�����ɻ,��XV:A��,!?A��Դ� ���&������r����ԛK���X�$+�r��!��m�@�8po��;@a9��V���n[e?��#������ʇ?�B6���M��J3��:�޸�w�7�w������B��,�����@{7�B���OjȤ����� �7��L��{bn$�է,�SaF�Al���,�,RNѽ3� ʢ�< ��͉]u`��G�1I��a���z.KԶ�ky%f�砤���t��7���LX�[$aw�R�Ik��GB��� ��q4�`���*�}S�^l�i|a��T:�Ss�H\m��B���KL��y�����8�c*Հ�Y�l��H�	���cY�aq֛�}1�\q��۷툚hx�X�]+���"�@�[.Z�$�3���mD��"���?R�%ی{�N�u��at���y�⾛t��?Z1�B܊B�Mi:g>��2�Bu<C
�b˲�����F�}T�HS���c��cd[��2E}�Ix�a��H��M×�0�(�U`����w"ht����h�㲪Fڍ!Uu�klHE�j/��/�ҼU3�=Љ� DZp�;4��> ��?�ܾ��	�N$�7)��� ��^��d�D.��	sW0]@n��6
�8(��R����e��� <�X=E��\�h�j��EWwދa���(K�I�G���Ҏ���_05�`5V��}��/��Ҿ��ju���p��a�ڕ�)��e� �e��[�ŧ��$
�A��ᆑ�"�؉3��6ı�[�P���j�}�i�=
��`]\��n���(J�U���vD���^�{᳋�n�����~�c�J�=j?�ή\���eBH�W�v՟P����^Pk~�v��J��h�w7�ج���v�����㒼�&�����E���f���⍊5�љy׻�Ӥܨ[�~�SM?d�ǿh�,Bl�gOX�	Ap�'�&%�G�O"�P����nE����=���� �K��2"a�G/�8.��j��8���l�F��?2,���3��;ٝ���h{��IK�{�g�x�
���{��h�����k���@�����OA)~��d���ͤg��s���q>G9ؚkdE��w����6^]�[�Ā����*l���3�Θ'�pxR<�lM���oA[>�_J����edn�C�ꋌtp�����H��@��|�@��&�5>:&�|�ו�[�����"����k9t�QID%�Wq��q�*}�Fc׃����q^� ��,�K�-�O`6��R g� �9%p)\��ئNT�ֺmeޖ�C�3��uA�����v�g�o^��%�2�'.�;����&�?��Y�7�hn���)��fZ���|F�s��T��PH+z�k��ċ�����儋�`�=�k��	^:w>�5��l����g_�l$G�P0u��	�y��1(o	�͍ ���������$��@�zl������'��V�c<�1�e6z������,��9��?TGfv?^i|��Y�hw�k;�Fl[��
|�i������\Ʌ���^p�vZ�5(۸��6d[�s%����j烶�☞ǯ�����L�K(�֞v����������lN��Zd�#��=m�p��L�S|�n8�	g� a++c�5�؋����1�.C�ސSE#^��V����)m-�x��-7�8��a��4����Y8B��+j���O�Q��PL��q{�pT��ݖ>�:��,�{oG2�8�"� ߢ��{7H���̓{*'@��S��C%���dbx�xP�櫸9���+C�ВS&��� ����*;���}�t��5o5o��sg���Ep��D�@��Z"��-Ǔ���c�#���U��p	�`���C]��jtX�^�ٴ^)gZ��\n��۠��2�����\X�|��bw�p���ƶ�����}���������^q���	��G��g5Tt;�(خ�ܾ�S{�[{tq�'Q���_E�x!{8����	�oQ��lx��7C�5x{��l�Av��G$mMDdo4`N�/��ԡ��o�g9A�|(�@���@SR��k����j@-/�kk�7�vA掐u]DiƱ����r����|�[=>�����xЌ�j���wV�������b-S��*��]���1�IR,1�1(��� 4Y��_�[P�j�}G��2�![A��L��
�Ɣ��/�Y0֭��E��s-w�plފ��ў��e��&��]�✸�2<�^}�"h�/�;d�x>�4I���#��{�ăM$;/jL�m�3n�-\����\ف��=L����r��%i�z˟U�ߙ��B�9�8��;M����^�b�%&�]$��۫�˗5]U=1C��r�h��N<�*~塇��t� ���>0�,P�h��*�m�o��Lj=���{��D�$�.��r7|yԂ)j	:����#pQ�Њ��&�.�o��"�e�׋b�{d^(�RU|t��Ⳡv�Ŷ��ا��O,��!�4TLO���T���/��Fh� �x�8/���>��Hp�KЊo�ݡ�1���n����D�9��6���c?� CR��?:����G0�9ZI��Wr�oP���Z��b���wLnϙr�m_�Z;�O��+��]/5�z�P����Jp��H>������nYv/��yܘG!Yj�n���?�v5�����P�ٿ���Y���V�y��T�p�ݽ0��X�=�	�pX�<B�<���7V�p^�������[X��@�ȸ%�&�QK���J��_L�0���f��GzsU&�n���y��Ih��n���c�y�������v�md�v�l��(խ�o_�X��!��ڌ���Н�}�*!�aS}|^���-��a���T�=n礁%v�󼲇��� [��I� �W��aթ3ε�XeE����k$��[0�̟LQyz�n��ߒκ�mN��~����!�)�=l�@�F6ț e��/���|�K"!���s1�2$V3K���d�m�Vf�f`�P;��V�!�#����cch߱�(��l|��?�B��S��k�GR��T弪Ry��g��m�X�q��_0K���}&�49Ό8J�Aod�����pC�-k����၁:V� �X�����AF XE���8ᖹ��f#�(r�zÌ.��؅ľt��F��^c���5��Ӟ{�_H�f��P#�3)[	������Hl�qQ;}���s��*`�����4�h�)�?�ЧnYy������q�5�9T<<�J�ؚql�UW$����
��R}��<�E��&��$��Y2Ȉe��'�o�E&;�Tf��O��fE���O_-������'K�B�08ܤ���IQ�SR��N��/�`9�� 3x��ۼ�E@��?G�X�±]��mQ�n�؍X���݊�XA�����<9X?q?�Ò�dU_fg�{��r�AtT����:}1�)L2Ձ��?�����NE&D���|��^6���f5�b������7$���cy3i�;�œ���r<�����sN���
J_�S۱ٞ0�∥��1P#���\��IY�u@�oa�NC��\D��I� nn睱��O����g�,g+��e6詾�حu�S_�����/f������6��6]�:?��.?'����o�,(}�ى��s|W��͖��0�UQ7.Ξ�ʜT�e�[�n\1�
����p�zP*Ĩ,x��T���":rs@����峙�+���^q�'4�t��{ǡ{P$6��q�v���Z���ߎ�R�F�Q�0Y�a�����8��7	�Nd�m/��7CJO�^vǪo��!3��ĭM��&�qA���`��#T����A�0�S[���F��6���>���Jt��			g��9R0�ښ����f�������CH��Hi����`�=8i�S�B��"�������Դ^'e��|{9Q��~Ym굾KnG�T�|�oo���g�{�mgR,}I9W�ľ#Mǳ:��3��x�N<����/��𜮻�/�_ &�(��#@�R,c�AZ��Y,.���g��yX�,f~<� �,w�^K�u[M�Y9q3�hpkp�J����h��a��%E^ ����"'�줚�%�$�´G�i����w	z6V�Ї�U\��:�9��J�.䒴���{�\��q$GAN�V����:������,�Ɉ�����&�$����ki��EE1���e��Y���d������=!�����k�KĤ/�܉�>m#�T�&XZJ'9(�;7����G�r��5]���:���NZ���ņ�_tt������z�+�78�4�4���԰zz{1qqъ�"���O+��{�:.++�c�m�Cg7K�'%�6�'+��.R�"���ז������*��Јw��/�ID��q8WVWO[Yi0N�.�SY������N=�����Ǯ������E��$ՙ��Bl��?�a��^���q�`�p/l;�����)��$� �Ä�TQ�2)#v��?lOOO<�Lܠ��2.�,�Q�}���@TO��}��H�x��%�^�]Ɓ�A���m?`g���U��CQ'&�##{�|O�1yz�+�mf~�r�����n������ީ���rN��CǷv-x�GK6�Y�C��@�Q_E4h����)�Z/���Vw�������mX�͇5Fݢԓ�gá�3�;��$�
������J�	�+�eH�?����⡠��[ �sW:�kT2wq	�a~{�����;�}}�����d�ݭ���1V�¾���t��ǘ��T��|�|�/�6��B�y��V����BR݄��?*Kϩ$syl�R����zؓ)�Я1i��f�tP��t�o���J�k����yy�R�./�}��[��y��rSA��g�D":�?~��Y[�C��q���%%�������#''�q-�|Q⤹�E��mc݂��u]��TINK��߿���Ѹ�Yc��SJv����555@���8�j�D�t��.��ٱN�ٰ���֮'���v��2gg0
�@���l�wU.޸`�����ߦ�B>���6����q��1;�����8�w�L�����G�w*t�?):�='7�����<z����H 揊�޹�|f�ƅ�\D(S3���ff�L�zuQ��h��c�+�2�B�̸4N|U��[ Uj6�1%�Ә[��Z�C����=NQ���6���ƅU���S.��< �?�k�ܥ�R�l�k�~��tff�p��ݠ74����G��m�֓�KG�xs�x*M�z�����i�9�f��^p@hs�O���C�`\�s�Gv���PNLLHW{{x�Sq@gg����m�u����6>�G�ӕ�3��z�3RQ�i'�~�9c-�S�t2���5�l�(z�͍����A�d�-0)�R�w�ζs�O��10`��[:Č�Q����;O������=j�u�������"B�5J�0F����U�E���斗��铌�|��_o�i~�%���<���C����� &B��/c �ȠىF^~GVV����~w9����T�L���uX�^�p��>�N�6��²����&o��{;��Cã�ţ��U��Y'''�Et��]Z���h���憻iwc#�*�%���0R1K]U���Ĥ��8�CgUUU]ؔȌiq��s��#X����uWIKs_B
�g����R�tBGF���-�Vf�{��q��, H��M%����2�
vv�������.��J�y�3��N	��m7 /%���Y������瓩�����U�#��/n�پ����[�dx���oED����&Nwu�RSS�}0���u���^�VQr��6�a9��p��{O`ʡA+l� T����q��#q���	+5#rw�\��'=h���떶67���vx�F�ץ�й����>�MX�������7q"�Mb����O�����6<���Ԑ����Y&8�%��x���.#*0���^�?�֣A�d��ajΗ*�b�:�c�k�
j��'i���YNi��Gd(`�b)�x�����(����|�..&�{X���{�?��ҩ���av�o�1��AE�3��n/<-i�����^Nz΁��[q�ᆢw��L��	�����d<z577Ҵ�j��J`�0�`(��忷tA���VoBґ���3q�3Ӽ�3�@�)�F���nK�t��D�@�E�����8�}Z(�:;� ��{xH�yׅ�5� ���Z�d�XG<�EZ�EAE-��x8|���6.9��ve}<@�|y�#�ܑz]{|�B��c�_x?#""�14{f�T:4뚚������2=�@񇧢7�9^���3Z^��؎��#2�zw)�g����6aFF����A�⍧,%����2R���~���;�wA��vrb�Q/��D�'���ښ�kө�!̓f,��tީU�i�A�����%�Jc�Hz�F�1���2T���7ὊWTV���W��ڃ�P�� Q�o;~��G	�	�{!!!
�*n�}BܨI9ʢ[&� ������=<�I�[��f]�۞fu���+��Q�R qO�l�XYYy����y�ԃ�� $ģ�
%�өo;��6V�J���b���<����!/~�Lb󣣣��Y��,DLL����ЍQ7���ߴs)Ee�S2�0
.\�yIIa���}��>���ɹ�-���,�^�?z{y|��V�i;���W��g�X�\��x�S��i��&���e���Ayj�YETV,V	^.�m���*u�Ƥ��ڱ*����=��['�ks뽮��T�����\m޸m��ٿw��N�<��Ej��g��F���#sNH��-�#�FD) ��O:?��U��PtQ�B���_�P���y8�����1)f�6��^��<��r�3�����'�b�Fަ��%"++ �g�%[�E�t��8CP4�LIۭ�0C�_��I�~hĈ������*?�fF[���W�
���\�af��;�t��n������G���C�q��?8��,5aއ�j����ʆ�R��W��=Ɍ�������A$�)Hz�sԻb�j�$e7cGA��ʴ�=?A�P8�T�����H��eӚQ�/�}�l����=�Y $-���wM����^�.�${^v�$���2��4BDK/ ���ƭċ�̃���*��+f����T�iL��p��I{�r��F�ʡ�@��l��/b�l尖E���
�_����z8+^��z���v����q��)�
iq 1/444>-)*�y�*��r��Цf`t5���9VW�޾:�ݖ�"~�b���xbU�	��і����W�����?������0��87�t� ��ʬ=Qs&�5�RPP�U�'7�u�����J�����C̉K��c$ߨ~(Q`#Q��g xl �����R�E��^�T��5�;�X�⽢�k�`�G���^�	���u���T?|��m{{�A�;3p�2�H^urNFFd�&%���i&���	�	,�m
�-0A�����[��:�_�Q��f��>�L��=��)���$�~�����5^{KZ�أ����1e��bPD9/��do��4l�<FH�pD!����b���(-��fO��^�;�A�>���Fx��y�@@.Ϟ��mn��^ݼ���{�����~�K����a枢r%/>V�|
�:6�sџ!�0�2��O=��L��ouuu�srоg�eK��?~(hpke��tGNÅS����+��b�c���
��ć��+`��9��RaaR)�~\�%xx*Jv��R�&G��Y���\2ldaS�O��Rr�l�����:o�����!�m�p_L5��]��><*���P ���b��o���ݖ�I�e�?|�( R(l�R�}�J�Ϥ�X��J��`tL���9��Ǐ��H���W׉�j]ƵVW�����e�y\[Mg�닯 0�i�1h:9�W��t9TD����t��?�'[�����X8�����5'�;������dyE%��rsG�W����9=�}����Č��-�,!������𩪪�A��K���[�k���5Tb��V~f�kH`&$�qP>�kttt[�vl	��<�M����|m��#`6/i~��������ָ2���n��o'�|��w8��k��T!H�������b�,��^�&dΏXri�.5/V
T�F$D�ԥ�?���,+�f,q`��EX�Qg^Rj���O�&��:\QT�Y������:ӽ݆S�|�#���: ���XXDW:Fx���
���@;��D�(�\^^Ҏ�� �O6Y�O��*�GIO7R
H[�lX��>>��;�S��v"���z"sp�Jh�Mω��H�a�(���琽�^2��r�O-�Lr�5þy�a�v�XMtB��/��Zݘ�A�j�g�m�XB���t]9�[ʆOF�b�*ggQ����Be��4��}|ؔ�ŵ�ѱ�����`��13S��۸v�:B����E��ƞ��c���oy(�q^�&;.���xQQP@�%=/2�������!=��l�;;�rN�M�q�h�ƮZ*��ߗ����J2pݟ� L�������NN�Mr���}X[�T���G@\P����)�ޔOM�fk�?.�O�q��E]v��JRF�����$�U,C3�S.qu��8ͤ���ދ�hs^f��/;��$���($?|7c�I�&O7���1U��t�}�q�«���/g7KOL`"�&���t�Bk��A�}�;�]Z�^�&c�@��|jLr.8y�&���������	��fK�eK37> G�C
�T�=K�����a���+���R]\\�厍)o-�׷ ��M�N~2:�8NHYH,-x��?-3�¶W,�?��V�D0|}ݰM��E���JBJ����w�&�o����=55����N~q��x�-'��8���hK\���e��iށw���-`M��V�-h��'	G롤�~j��P��,|�JJu���Q�wo�;�s��Y�¶��j0uH���-��1�L�D��^]]=s�kr��-�795�C��-d�����n���0�}�FoO��	�S�UJ]�Ow[d��_�'�3��K"M7G�9���gRc~@�O�{�}q\o�df"��q�[�D+ێ?&������KL�8<f�/�4Z���9��/��,��,�5�>3GG���N02k���=kkk�6L� @��+���lH��l�� �!*�,DC+�� 7��ҚP��4:OK��y]����$x=�?/�;��45���<�����[?ܳp�^���TK���i,����"�?2����rrGG�\hXXBnfX�_k�"��͋�3�	��6�. �+;	`�^���+z	�=�"!#��#%�C�ُ��<0�ϸ��~�7J�����NHR�I6n���X˝�5j���(�+V�ޞ�_�?>+��b}w,����\�ݗü ��Ή8�;�t�|q���}�f��	�͚s�����/��WY�o��^ E�\p_�a�C���ݏ~�	Qz����E��M��M���W D�|���ح���o5�=��JPM��B�ioo����}�V��l�,��^� )�F��q#�޶޵�7��m)��c3�m�����f�����h����g����m&��Do9�$qV:�*����`l�P�8Z����(�x��}�͍�n��ǔ���H���ך JRRm�������q���=v,d;�Z[[�ѽ��a)�!��`~�2qܷ "�D�J�ݺ�8���D���0&B��${G�r}C����*���Z�{R23����_g�J2S�����mR�a��=b�B���J	[ݬ�� ���))L��|^���|��=#CπK���=.�0}���K����!�8	������9���F��������
�F�%%��͞�H�ډ�]*�>����9�aZJ&���)'�.	2v^�7��2q����X�B`��������*���(�j&Q�z&j��> �%%e�{:|C��x�����2�52�>e��n�{�����>x��e)9��ޣ��6܉,��G���I'����o���qd��a�BB1'՝�:6� �����5.� /��c��G�- z�hMT�m�99�l�\(�nfV֗6���V����`��[�8&�3G�k���"0�0����	�Q���-	~i��g��IQY�����&�N����||V�I����HEE%95�R��u~����㸫�n;I��'��%�8��w�ei����%!!!��}[�#�x��  
����eff&<"�[^���3����[pc?ձve_�R���j�!y�F��S+c�0yn5[�a644�R���	��g�F�5o���%7k�@�Ji1�)W�w�'�������]]]�����yE�r�ôQj��D����$0�bN�z]�앶6i@�/�@�1���$[v��|�i�x$1yrb������/�J:�CtmvQz`���F;��G���~"�&(2�o,��ӥ�v����$"��,��2pn��Lʕ{p��<W������WP�Wò���S=W��pi����Ftq		9���~X�)5�}Z�_����wK�nj,�����O��h1�j�ד��q���^*B��=�EV3�����)���,,D�-뢠�����29�0 ��O���-�&����x�ӢV�O�D<���.o&2	i��ĕ\���ka�Bx�wQ8���B)���ZN�H$X��p�-��q�����L�*�;��3�/`���̈��O����]����@�?uM&����+���K�W���w �:~�4�|�C�(���{�����Qy&��`oo<W&�y��l��CL����꽁�˴xPѫ�\{8�h;ی��rR__Oǔ���#�#w���_铌lm��V�4�Z���u5*ϐB����ݿ!v~'�q���die(� 7�q� ��x �E��A��͵����`yP�y9�1ȇq/I��ﾨ�_�R�����{g��,���<��CGY��JQ�:^����n�qa�|���JՁhL�n}M�� }b���!�=7��tSVfig7 ��g]�.�ʎ��I��e�����A�B�o
h[��}~��ebd�!����OH
�:rp�Q< �:��W��I��<G`���|0�cy���'��{y��;��Wѝ�7@J�~�f
����������Ⅸ�a�"� cJ�;V�t���|Ej�
��%)$�$+�8b�7Z@5w���������9ơ>W����(µ�� d,h觻Р�\��������_7��;��w�w���u�3��Z��m����~6�+�@�>x�/���_�1�R�S���"4��Ma�Y�$Z8�WՀ�(9�fE����!e����l�i���Tgj��ǩD�N�z��v!�o��m'������X8�
#�-�I'��tr������>h����+i�+'��@gq�o~��į�w��{�T� �n.����&��ާh*��7R!$ґH0����s���4@�ۘ.S�E^����;�SD�|�sc�uR�ow{y+��s����8���	W����W!XXX&��Np��B^�g��oܶ6��ᓇ���Ƃ����t໑�"T)(l��Ծ�y5���7W�#����~��:���0�O��f�
��������粐��WIXR\\P�~��l������~��ЯHN�\9D<_��8^HN);@h���Ӆ�d��Է�e���m�da�:�r��L�Y��ڿ��bD�SMU���'��E]�%=?�V����Eε�����ͽ(ToX��������:��	����ɖw�n999bѼ��FN�H;�Y
��0b��v�,�Q��Q��!��蕙�3���8,����W����q{>�d�#Bf����C�k�Q/��S!����"+7���LNn��va.T��1	���V31��������-��g$�;���o�u���V�,MO�Wgj�'&��k�>�
��W�"VA���̕�"�k�'���� ��u�7��~x����%6�!a��ɓ��]*Kv�N���b�͙[X8n�P�]��%�����{�����)pU�no�*)����z����[i����b ���-�/���-�����X��8�G�#�@�i:�e�k5� �i��"��\r_�ig�Q�D�􉹠�@�#.*�w��(��t[e��0�
�	p�43j,Vyr���$T{%"y;閉����kN���L�̍���Sc�rUu�1��3���� 8�>'a. 
�N�|fs{�0�߸�|('Omim��rVY`���v�/o�}αaЯ_-,��R��[a���BQ�$}%�~^K�*ԓ�C2To����! >9ك�H�^�	���J#"��i�0�g�����$$\�ڀ�~�l���$������G �tm����������5#��?��쟞�}`��`D���|��U�)�U���޽��w���������`�����BK����$�kAL^s6~������	cB�m6M�������ӗ�1�����8 &^��A$̤�:U�D��N��Wy#k���׾u�V#��N)��gZՊ��hD�utl���V�������f�P����a�����;Q�ps`�,����`Ak`bd�����mB�:���V-U�Q�g^^��C%Z\�v�b~���/M��)o("1f�p�0�Ђ]蝙�)f�����I���_�t�P���s�%)1��ʗD2Ҽ6o��(��4i�(S���vu�}��w��ґ>4-��
��S������Q�>������ �*�2����p��[���ĵ��C����jT�M�P��6����mp?sre4'��%�}G3��U�?)���#���u7W�(�:8��l=1c�b>���_��&�p`0Htj7�Y������OH(,>_Ke��b�� !K�����U(S'�?O�4QEM���)�^�u%`��u���W%��\x?���bF*EZ�4L�`�UYY�&$���U�#�k����64�����p���|%5��'J!��D�+0-G-3c D+׵�=��9@���m�022�57lm����T�O�`�d�z]�Ł��wCoQ��y��}�\����'9��K��VW��,
h�k�)�E���OϤ���4��5?P��~w6@��U���������i�
vGϬ���N�Iփ���M:3�O�̹ffE�gߝ����������/�lM�א�^����h�2�fkP<�d	OA��/wWd�/��JJZW��\m����-������]�d����#?������%�M-J�������c444�|�e��!@���I0��N<�h�(��fh6=��D�D���X`����y�!yDO�2jN�	��+{����f��0'd��k�$l�~S+�oUR˴��ի��7f����m����;!-�F�AK�[�H�E_���
�QY��4Xÿ|�v��}�7���"k~�FK����J����:��3}��+�p Zd�A��TGH@*��/�`���lR��̲I�hǵ���eap`�B!�s2�|���=���{y�|�xv}]/X�M	����>��z雩�!�-pI�!m�C�ՁX�[Z|�d�r�E@B���%.R�J}��<y�t���Q�����DMb5��:��ښ������
b�ތ��?�Vc��z=�c`f��{��{L�͖��Q���t�Q�ʞ��58(w�S @���{�)v�U��>���������G�	AEE�۞Z�!,�_\ <7_�'6_����?�?�I;[�@'ԝ:p��v?���7t256�Jy�LN�(�i���X�:H�Yi�����M>��IPkH������`9ͬͅ-g�^���<zIr� ����k�1��i��}�յN�{=�`�;;��*\-���/��V�Դ�1���ɻ[�[Sb,+w����g6�@����pVj��e����C��ӹ?������WA��_�8��Kk�?OD�6 *;�!V1��V���։�L;n@Tb5/k����ָ�L�<�~��>�vQ�/����F����vvv��'#���L�X��c���9���#������i����6m#�؎̎�m�Ě־p���QXM�D�YSG����(d�
p=}M�@�k�d�OϷ��������k5e���ǟ���Q8�rpL@� �e�/U���f���_e`���AZ�vcqy�G�5��k�ze���:}fM����n\�V����6��W��1�j��"�0�p����������%A{{��Ѿ�������������ە0!o������i,k7�n�����*"-�����{l\#��`�IV	Q�dF%����m�1ו����V�X�����ؘ2�\g:�D����������J��()e!O�
/�Dkū�fl��v�$7����*�����*K+���w�׋���P��(Yx�rE����&i���%\~.L��س��� (;)�qI�O���\M���.'����P��՞���nC��nF�H������).���1�t���)�F�Y�ʾEW���S{�JQ� E��fg=ܨ�Ycͺ dQmΧ�1p1�_U��?:�B òD�ܱ�y���~�,u�1���9A�H#��(?�`�}���F~V`;����#)Xe��w��>� �vYW���J���hj?	E<���E�C���z�w?\���JTu?���� *��U�$d� G3�&>�c>C�o&_Z䫲Ch�5���U*{��\N�ѿ��3)
��m��<�W�K�5p
R`<��d��5��y�5����g��0Y�^z�͖����]�����-*
��[h�o���M�x��z�5����n�ٚ�yy�1�9%q�WR��0�����|��"���6������f3glhh蠡Ɉ���Y0��k��]� U��N�:�P$��Qe�~�n �����{GD��`*��3��{�:�T--.6�m5���=XGaO8�k�ú٬� Iѫ�V�$�
&����y���O�Ԧ&�6X2�b� K����C#��?w�씂v�p{@�ܘ*s�`���i�/m����v��*�^qykk�V���|�����`f�:��\ms�aI9�ϼ�I���DƏ�bʱ��Ĺǒ��<?��SRR%���0|��[rJ��f�����`pH��G�=W�;Ч�&a�Ϙ�J�t��H;ǟ]���Y��i�W�����6��N���^V_��~��|:u��&�\inl4�G��E��o�ǈ�g[��l�6�
�OO�����>�覣g�?�|��ګ={��[�#yy?fd��uPRӄP.���I��K����Tp��B��g:����B:���-�"��6l�;���M()�����zDi��:]8���3)�1�зN���r5�����k��+���n��ֆ�>�7�F���V��]j�di�Z0e��ʝ0�c%��9p����z[�+*v���� ��O����.7�>,�r ��*�t�N�u߿�
�Ce��ʹA��T���^��K�2W�������2�ߓ�3:��.[�r�������}���P�L������"(�fd�i}�z�U�R����������ԡӇ�����ϝ]�脴�k�\"���$�c0�=f޴�����q�K �
sr<��n�/>'Ci���Z�^jk��?�Q����ǌU��;p��{���#���'��@�ӿB��:�%�,Qy�6��1\�?�����ډ��=� K
3'�#�٭lE�<��S͗�\:c�ָf�����ɬ�z���D����FZU��
���;H��-�޷F{�_Qt(y�yc;����g))���gdg#���G��=t.~&��|@
C'�8�! �}V�.��G��w-���A�5#١<�������xg	��2�}�O��B<k��I�89��]  nZ�ѥ���ɈZ�o���h�F����u�:s#�" "�ն�YnV�O��.�~66�̀؃�?2e��� $"<[,�VMd�=�]���~��ix��.���$#���E��UHR�]���I��b���;��)��'R�$%#
�e����͜�1%����^��Ԧ�«��@q���~�_}����f������_@}�ۍ(��(�t�
���k�0�QX����ck�ek�QvV֖�4�'��µy�,�������ghgX\�� ����ތ���ά�W�u�\�zx|�9����~M�Z���;�)�@��~A�4<.n��&����ֲ+�	��4ꗡN8�z��NC���S�ݎs��M�m�� �Iڟ�}��Qk����D�!!g����������E�ړ0�������[Fe�um�
�Hwwwwww�tw��"� ��tw��4HwH�t*�{]z?���1��w��������s�k�y��q¦��2=2�̾��h��!#�;a���g��Iֲ6�����M25;�R1�B4O١��TT4�U�w��I�"�Y��,���s9�ڻ�980"�ϾT�/IMܰ�����#�o��P�Zpk+_Y�Z$&}|zVد��tòIk*����,�FR!!��n�&�������T��go��6����#w:^ih<wm6`�<^E��0���T����-*.N�ThZ}�B�0�ۮ�.Y͢�ʪ�_��<�z�KJqg���ThX�e@a�����6�Y.��P���Y7��l�|����(�og #R��0w\[�� ��+���P`+4�5˴q�$������Z��^?܇"�5�		�nv�]\^�s�&ǊJHϒ�=���u1A���=�i��*��A�|�oFɋ�0HUh��{㠕̔o���FHD�R��=�(r��� ��	��&a`�y����K�h�G��� �B�)B�Pv�LnT._�ixx����~��;H���S�֒Gtt�����=D)~:A��O	��Vc"�B��`��j�~�o�q��-�z{Z�R(��O�|Y��0��룿�#�L�ng/���:����rrH�7�x1�a����~S�������> ߈ ����:��(��Md����@�Pk2�l�Q{d�W9	)�4lxxdqss���ca��KAAU5:j�*p�LCi�Z��--�������eʘ�V��?y��$y�"1k�bg����l��߼p��/�����p����}m�$��� �����W�?�{���w���ҁ��^�|/H��䉎�r�)�v�Q2=b���g.�01y9XZ��Gu� ���3
��v''����6-�}���͂S�L?��q22�ޜ
�g@doBJ�u�Ҡi$��̬������Q���R;�k����%x����n�"���s�*�	[*'��(+d���zຯ�U�w�Q����r-�	�7c�At����d�!]
��ϯoo�Tc=�p��$���L^\p�ҕA��8��R���!3,��Y�%�k5�zF����Y�`I�����>�X�䫝y$څ�������%k9��4��@=����M�/����*���픺i擴c5`���ŝPRbϱ�'_U�i���%3hu*=���#�g��O/@d�^o�@z�2@�Gy3r��h�ʗ'ߢ�L�rv��Ē^�y'��:Gs������l�X_j�8eE��(bEE�n�)Y�j!u&���JL[�A��+&�5H�N����Z����ԧV�n���W�Q�z�О@�f>3�=!ofgaa��_]5r�t'�������)?b(�5!����>SU�	��FH<�ۄ�ė�1%TD��dd2!���!K�L)Kh��	�� �ϳ�T�Tv�F�slm����CbK��������EXyڻc^@�o]��33�Ggf0���ߎߎX��������.����Æ������&7dn�T*E�paY|���l���#�|�e�hcP#!3���Q[���$1�BZzzO:P@aZLh###٥�p�eZ�4x����q3�&!]�n�Y�ed`��c�_�7ڦ���舘��3�p@Ɯh�j�)��Y�Z0�d��y�S;D�xuw�q�5°��"��G�d݄� ������F.k����.����*�x!�y`�4�f����[G�"d�)�Rn77�skre%
`�nH��v�"��Ʊ	��BJ?�F����T�&,1"$"&����#R�A��)\��^�>��yVV��Μ�%P��+�SK�C�p�)6B+�����C�PvI;DD�0��Omǈ>?�uY�;s��ߠ�����m硳Y}��9��o�{a�F3D���e(TJ5RL�xiI���
��9��R�t� U4���B��k���05�/�F˜T���,ϩӡ�}�������ݬ���M��pS��V	����Gd����O,"��]uwC�Ce
���ŋ�'V�҇-��~k nk���\u��fD��(�����ȇ䐱X�2%_�jee��a9Ttt3gH|mf~�����-�X&���3��}��I�����ɸ��3��v���>�I8��zZ��a�e#ߏ���	�f�<6��L��j����~tj#a^+E��'m�.%%51���m^�,���L�8����đ�x���p���F$!���аB�v�mk)\@��.�X��I�5aүq������إ��n�&��)f��7�����ĀDb�3����|ɗ�a��������V������[\�i��>��e��PY���?Y��#V���8�����v˟�a�5 �<T�h�PBp�Qլ�y��K��r�ߵ�C���a��	��
�T�XS���dč�(��^?-=!�c���//@�[�|YY[Rō��}!PD�@��+t��MV�Ww؇���b��s�x��?S�
�9�~��{w�X�@m������[���0��'�����4��T�����Bj_t�m?/U�33�>e���LO���`������������#��Sqa�HUK
(5	���XY�z꿄!Q��h$����la~n��������q���	���-�JE%%1#2��u����^:e2�)?�ݯ��	����i�Qױ�PA���'����3ǩW�`�S�[9��ķ�;��Rff��#6���tC��!5�y��He�߽;�$�����2��g�χ$�*)����h�2WwͿz�8�EAI���`�I\=���ď����(����}�Y2���%J�c��^� ��ar����w���cUh{g'w �crb�O��BM1J��E���д{�(��F+j�N��5�z�l��,!Rٕ���-��^|{.�o^G_��Lj#<Y����\!��dk����qL��:8D
jj��I.��jͲ41y���rz�,T�5�(�5�j�c��ؘ�B�%^j��g��w�+��i"V�i����r�s������z'݉D���{M��◨��^�C����bc��I������Ѿ����˂Y[��afR��]��e2�g��̿��9! ���P���n���/�z|�VE)f���3!�27���/±_a�4����%��}�)�V��g�F��6[�)��i�鵛g�P&s�5����,�G�)��g,t�hh��b��!m���$	2�6����Υc�S�O���������XJB.��Z$.]�".���}\"�)��4rq��Έ��*�-���u5@Y� �.k�fV�,U�0����L�h���.�ߐ�P1TZ�ښHY>��5��/jֳa<0��}���F�w����j��b���3 ���^%����d�p�ڞu?d}���%/?���p�C����)�D�s���m��q����f���t�}��GA\�WЂ�V��a��jbb)qO[(d���֮�e�!ȁ1�xiDBa�>?uzvpӏ̯�~��Ջ���-ſ�mN[���f
�ԟ�OT��-O�'q�bϕ��n@�t4��1~�h��ө�l�\�UW�9�W��!��+�?V�|ݎ�6)	#o�<--MEM�~^j("�eFyI�ͯÍ�~r������nn�L�:���!A�れ�o�4Ȯ����G?�ݯ�Gۦ���3	���>�OpXnn�)�z`�h��E:�S����� �����10a^�
,j�9 ��������;2RO��*�2E�1�|�(k�ŪRد��b�,,�Emm]��9��C�y����>���	3�<B�K�{k�:�\dD� )�D=kq���W*�j�e%%����w0����w��6L�=��ԣw[SĚ*��� ݞ��v:��G�Y������m��Q���y��<�v�xA�wA^�H�a�_� LZe�l�8�EX��ֹB�:��u�QD�퇭C�Yl��*���qL������*�q��^=#����2?��͏��Q�wY.�X�:b�$�����x�d�Ų�m�R�����w�&l,��G�m���X.{`�p�p�3]c6������Z������t�������_�"���������mξ��ێr~�twX����I��(+s7sy�,������Heg��gߍ��[.��XǷ���ل���ܾ;����<��6ʥ� �*2�H�b�Q��b ���?]��;N�������U\Y*��h��� �(/���h����� #)�

��935��
�I9�fff�E� �e�Ѥp�X������ђ^��E_ѵqa����+�7� �H%F$\pg�%$u	��W�h%��MK2gsI-�0jǓ+x_2����q�r]�[5b�������r�`��*��
;��1���i����2,͞߿b�����ӕ����)i�}]����3
8���d����yL�b�V_p�����rq���7{5�{8_��D��	U��K(hh��Ʌ��2�
B�=og�o��>?d%3K��i��Cj�lVRü�Ӓ2��be%�����v� ���{.���-,.���7(�d]���]�G��_ގؿ���wX_iPy020d�Ԡ~����M�>P�|����Ӛ��^�fo�А���V*�گ��sB߿�U�<�����E�<�b����!-+i�^3,]A$�<6n)s+����V�P�?��g��]i*�v `|C�&�|�6��8Z�����3b
�g�'D��!���>c������Jg�I�A����Y 2 �,�؜S����5�|<ᣃ�'U&#e~uqA����o�)l���(6!��jw����h����cMY�|5��SB67��Fl�:e�����C��߱������flg�&x���ó�k�nη\��I��C���|yB��h9�Ь���[R�P2��
y�Oq>�Z�����6�6��LV�=��h�捥��۲>�ь%N&#�4�
EH���$��ן�Z'������F�4s�
4Q�7��[&�Ƅ�;N����^��@Z���R��;%I�����f��g��<�'!��(40���|c��,�o�^��rk�$Q��v�9����}�4��IkN�x��N����������u�b�N���O�y��E٭��'&��n1e�ǣ���J@`�\QՄ��۲��S��Y&i�I9']A}������BF�j#��_u�v���N�7g��'Q�؛UԨ�����Zg���?��=%~288�Ң�7I"�L���!�.�x���'�!�3jCCC2���˿��2��8�8��q��сK����&%�i�������B�����8�$p�7M4geeu^6�j`�ᆛ�t�gw<+Lo%"�i�R �i(4���s�3���f3�c�ّH�}_ߒ̄��7�1�6���-v�hb.�%�OvU-R�FJK;�M�|�~k�4�ܳ��\�ʘ�R�η\�bM��3bZ����Ϧ���+b��c�_�8���ȃ ��{IHLLRԳ�w���͕�� i�>[@����c�2�I}��K�x��ᦗ:3�����0�hkg��G6�L�M��J
«�sʹ��t�O1���GD^��o�a%������3����� t����}�-�(�%Y�ߥ��W'��AA�U�.^XT�j���իW�_��f��l�jw����^B~��^�k❀$�������!E�)�`SK�ł�YP-�Bn�X�	XW���hN���?���$s�����F��k�2rik�s+ww���8��H<�	�����i:o_߃"ݾ^�?i�f;;�g���&&�J�w݀�)M� /*TL�OL��%�t�I�rN����Ͳ6���4���ȧ���Em���0FLL8��Ko̤�tƗLZ�}@Ȥ�5?pӢZ��(+,�J���6�=A(-+C���Q�
��-��۸���(cG5�����;������6�S������(�d9ˑ����l�����x+/���Y[�c�4ݙ��.{G��n]�"���g��3��w������@2��g�)��5[c#��� ܆K�MqJ�n������>��I|o{���7�]\��<�9�L���71��	
ƅ�mN$W_}���)Y�|�l''�JR����������7O�H����~|k����� �޴d�o�7ۨuh:��u�v����jɶL��)ͺq��3��=��iFt�����?_�'n�v�����B��J��n�GtB
��*�ˡ$�\���j4�;��};@�M������Ϻ~���Ç8�����RM��)�$|}VY�7�#3s{R]
N�������"$�,<<)�X�o�%.�a�BI�ȓ���˝Q�p_�'Zt�[v�A����o�dn^�KC�|�,u�;*XĂ�<�K���;���Σ��N�-��K���v&���ZZ�x���6Z��Y?w�lH��mmm㓓C�׍���͎6�m�����9����c����Ot�ޗ�����λ�b�A@����t����[�(�?^HI�4���|/���=��xc}]��L����E�&�|'���Sh<�f��B%�.B�Fn�ހ�
W�%>�b��7��b[�/�#N�z���Ғy�Ч�7�I�kl�&r`�Pb�c��p�RE&�M�)1-bLJ�@��&G͟����!��
���V��H�S_[+��;vL��n9]<~���ZFY>�!&f�Ti�a9���O=��*_����D�]p��T������a�p	K�"��!��m��(kjxy#zu�6���k��d �0b���l�Nb�0ɓ|4�
;;����5*��I��r��D��v�E���>#�~�TFN)���`f+2*3���Q�0�R�~uMMȰ3v� /?)	�]��b�R(�t8xlƤfY�����µ�+��{���)%%$GN.S�	�G, ����hs�𐕇�+�p핐̫�UJ*-z�??gʗ�T����r�;2�������d�C��ܜ2�a�a"���+`��/a_�L �<B_jzjc됼!O^y�����^�����yxl*?��6��oYi�������hACx���xICx���j&:��B�ß:��+)��I�t��ݭ�4���
o�;;�߫��S��*����b�5)��oav���q��蝉�,,l~	ܦ3���~���~�푝���F�÷�{�֏�S++1GG�˶�I����g�Mt;I�[,,,���涔��L�?������x��ǈ�G�����CE��n��S%�tEC�ds���m�h��q3@:�#"��,V2��.0܈��Oiw01ӭ��LD�:������~�g/4��=�qpg��-Ю��Ɂ*�˘A����C���ͰLN�g/�J������	�y_F����pX�$���;���7���h�}���>h/#�m*�/���"����YH@����s�������p�~�j�;��υ��^5>�T|�*�	��i#C�)�(���֎1��9p,7��]�4��C�����;%PF�T�3�r[���\���mc!,0�>y����?o�V:��{�j�
(I<=9q4����˃~x��6N���t���,�T��J}��/���R�R���Ж_�J(cbb�T6b�B��ېQyN#A�&�׃����_��[;8̪��N�9Pr��LM��S)��»�qX��IF'0N-ME"FD�$��%�V��������q���3�"�����!?�Ώq�=�<��67�F��o8XX<��֮P��ʎ!����h:���*�0�5�/.�'��#K���-2� ���n����&U�p�g�m�����1��*}�*�����~~y����d~b<zzz�)\���5:)�^L����M�^�YJ�9����o��s�ٳ98yzz�c�m\{Bur��	u1��dll��� ��ߦs;��P��`����&fd��9�̛i"_ز�ʄ��:ͦ� 	Ȥ��x��2�%ҥZ\Cu�pH	YY�vּ ���ŝ�ԑ��碠ڼ�]Q�ٯ �'هGQ�����a���1I^E%�u155U&Zy"J����Ɇ�/_yEE�ct6��M�o�>��Nu��e�Հ�D�n������*#�K?���2\�//�������o�tT�.��_����e�&�L����(Y�(1]n�}.Y��BDU��h~֋�6�"6eR�뚡�v^^�.�/ĺ�#���������+y�e_#�$$�r����ސ}�L�~SYW��̷V8��r�S����߸�=<@L����Iz���}�E��^Q��C���Ɨ�\e(h�4�t����4̀�,��W���++U�S�_�O�
'	���D!"�M�Uc�K SRb��4/f�c?u$	H��,�����-�\Q8S9|\�N�[���A���3v�k���v\q�	��#..��~8_y�$�����կ�e}MM��9I۶�?����c^u��~�GJS'��x���c���(����zt�����<D��s��剋O����c;��A�y�|��a �O���sp�	)�O�b�{G[�h%�!J�--��P��>��������ӪĎ�\�HQ�\#i&=���bp)�1�\֥)�6D!?w��N�ET�8{�ޛ�_<ݔ�KD��G�5���	��v�r���>P:��l����bM��.����*���Q#��tZ��Qߝ�:�����RPQܑ����rU�>2N�#M��6�ѫ������00H�+ �z�5MM�m��J|)��٪6��Z+�nI�W�5nt�"~=���^�:�*4_��GE�����^��k�b���
��8�[��+�6`��jpSTD^�$	Я%�-���� Q��V`�T?~��^����AE����`�`��@��P�S�	��RWW��'A��QH�p{��T��"&%�\���&>w��)�b_ ��������NZ��W�=�#5�%d#@l�G�� ���\�e��f�(�� 4>}x������$'8pw�?V�ё)-=�#��ǯ_�jrl���7��>�}����������$�S��������(~������A���њ�Vff�����Y��R��Tq�t,7�� w�mT<`	��`i�Sj�R9z�'��ZZd��ؤPO�>͘����m*�K����^U��6{A��\���	~�21��)-��u�$��C*2�RS]=(��Ö���Μ�b����Q`gHW'+⢁'J�S0\���ss� ��{ڇ?�4>;;K
V�cb��9�_Z~��j`��Yw�K����� ��Ii_�I��r��\Ձg�x����ږ@���1N,�
!���:Q�f�/�ݕ3X����m=U�����@Ǡ�&��Xx{uj6py|�ӹ�7�o�W��%� �n��KoŒ�2��ڞ�����(lk#�LP-.-�26/� m��{���h��J�ݬ�\�]os���pp%]`%W�~<�7O[V)�w�g��c���9�Ҟ�TC<��IC�%%���@ 0?Z��]���;ri�n�zj*,!,;;{� ?��;c��R�sD����^�:���X�|��3F�¶O�9��I�8�Ϙ�N�VT`�I�Ꮦ:����S��i����Ԟ�S5 �b	�3;Y��⇹����	eC״i�.��&�nO����}d�+-�#}�Rcg�
�T]�B���5��K���G�d)���������-��F�"��) H��lyD�Hc�V�t��+�FԺ�N� �T��O���T��������_����.�+D�*��o�;�=�PXM�a��u����İ7�J��	��Ȅ|�MM{�.I����N��yb�ُ�%dj 4�p9
v���
 |�{�(|m��{�:S%rrr�T$|tS���0�I�}=ؖ���88N���y:0��4C��'Q\Fv��"�p<�3d����HnV��r�7��NW�vӝ��E%��2!�ߜ"Qѩ�]��N��(@�dd1�GK�]����^�ŕ76b��� ��C��◊����U���vK�B���k^��QS�ws�]�]�(b7��f|�p�a���ي���5�3Dt��RJ�<7�����V����#^��D����)�����և��!�ԳP�=�E�����1�_�J��C �AM��ǀ	�^��wD���h��c�4��c��<G���Ev9MM�cj��B��ΟQ>�Ǒ	n�n?�� ��DA''Sy�ݢ�~r%�o" �9�����XCC#�Nph�a�����(�@�#�65I���-/���]�K]�9���!��g������b�2�.Z�wD+**xnvU����f�Y=�u��z��jRԇ����
Iww���!AJJJ:�w$������z4���/�#��=���~]�@u�����;����P�5.ݛ�����]Q��f��L֟���F�T�l,C�"dP���MWwV,_���@o�HB]�AD�48�_Z���[��ᅑ,�;�) Y�P��n{�M헢�|�.���?=������p~%�x��&�b�+�hi��֚��*-��E%@�Hz{����(�e���ٓ�p�6�����o'�����R������a*ŧļ���S;���$������� ����ڬKY������¯N�4��q��~���8\>��C.��G���q?v��?	�G�����~���?~��kk���'*]��/Sm4�0�d�i������N.,��t�f+�m����+Sx�vF��d��)�ǧ�gg���^î��4juz��q���9����o޼IM����
�m������� ��:9-F
<�'�h��|u/!�_^^f����:��I��V[F�.d��ߥngV������%9�2�0���|DF�@HO�^1M������Lp�.�*hXXX�q5u!"$"Jc����<b+BmV�� �ARZ���X$@���D<<8ar6����.��ӿ�CA"{�m�)��N!�����Nx��"�;�B~eH���[rZJݣ�<���/�o^�L� ���RX���)%O��K��a=]e��ԕ��V��,}!r0�k?to_YA�c��i�&&��yfB��-��!KJފ���u��a߭�Z��t��h-#,D��O��I��r���?\G��� B�C��ov���8�Љ��v�۷"itS���5��lk�� yu�1?k���s"��I�:�������M�yrffe���0��i���F��jk�Sj�\ �jg~��9	��Kց�鄌��ȃ��H�f�����J��
b\�:���z>W�t�02p#0PD�����y��E�T� #��iQ��� ��BZp�;��6uq�.'`�2J�bRd�v�3��:�*��%���`�j%t����Y�X�3E��]c2���Z�M���mu�p~���b)�Lm����X!:�����5�8��0�_e��`'8S��G�-����Y��m�"K��,�=1�|��`�oG?55���xg>���6�SV�Oޚ�I[[:`�8�Vk��ƀ&�=�&��Ѕe�n
<I.�f�%��qߢTI?�}�陟OA~�W�(��������!a�y��n�où���L�RgQ>����~������8=�t�~}�9�cr;��;��:�4�C�Mݐ'����Q�NX�l� NOaq��5�0�6җbl��g�q��V����d�3.��s��՛ig���㭠��DV�O<�@;y�`���@4��
��3FffiS?�ζ�����`�A���WL���K̭��̖đM�kXXX�~.<��4��4�7�Q#�����KLL1�g�&�-yEy3<�������]�t�,&&Ff)>�����-������
�|�:�����|�
²N�c�Bl�@�V��ڡv�w; F�>	�����
�*S��'c+ӌW�
�{����п�Z�Y�>שq�i`�p#?��b�a����Ib��xp��0p�g(KN��"�q�:U�T��':�LL���I2�}<�iZ����3���1k����l���8���G����+D��,?q��>;�&�*�x��LBDH��E�I��
A�#��p�rdU��H�I����ڊ:.$�:�})K�AywuXՀ�z���Lb�_�������m����t���vvv@�KQZ�p!>>��W9�{rۏv�����d��ۯ� ���sW�M���VY�t�� �3� �I�vw�QPS��k%>'�V B.�+������P��y.�4���E��� j�v��da:t5����C �(����"9������.��Bo�� �;���2��D�O����j+f����6RRRN֍.A����M�ֺSkB��˓`�)d\㾯�j�p��R��N���SLkt��~�$E�`ӷ3��\p��|�5��(�Ե�� +���06_��{���A��-2���w��➫Eo��Xٳ��'
.gMk�f���]h�-�X�^Etp���w�/Z����kӱ��Yhƨ���_��Y1�������{��{mh��a.���J�@������R�g> {ɅXEva��~M�;��Q���Y��s��β2xb�kR�sC�9�p��QQh~�(n�4���ʊ���sb���Cxtdp��Z~V�v������8%��\%jz�}6��}�i���������FG��$p�߱_�ߞv̫����l�U��(ʊjZ$�@O��SQA�u[���ީ�p���/W�d~_���B��v�+�Ht�h j��?��칰���-6����`z�Q8���Cj���#Vĉ������n	�
ۖ�2��b������=o�v��w�����[\v>�|4
��$��;'[)'������K�>������xlf���ǌ?��
 ���%
���P11)w�Ea'�O 	`�@�Z�t�;�C����݇}����xs�y��������o�D��}�����eЁ�]�����=��T��Iu�q_Za�
�i&i���v�%QGtv
�IJu3��=!�q~���7%˓�^j)��ܾ�[�ý����5���Λ�5�	|�����0s�׷��
���6���n�Ta�J.u�S��Aq�����S),�`��MF����ޗ����\F�F���l��o��!,WH?��D���KH��@FZT�S���M�1;:B\���l��"�6��)�1(��"e%%�b~���cPL�/G�?<�5;+��ȍNM��D��-����K��s�Ga1w��[��c�'�9�Ε��n�-�:�.������̮�X�B�ʊz��� �2���o
�k�)L,,2q����sK� ��WV#�P�l�����������zf���*rR!��`E]�4@e	#�7��M��X���
�����ϕz�A$���(�He�& Hx�~K��������C��%eˎ�'��/���Z�ՃW�u��>�\�����S������⢉�!!d��GG�a�~�yo.����_�� <������%��f�)��ѿG�^�*�_B�N�?�j1�:����/�(M|-���P����l��o�o�i�=���^�ݝ  �Cy�����$��>"LOD^��}�����t�t����;O��ƍ4�؝��98<&B�%[4��0�hpxTR�}��^�7}mml666cSS��-��2
��ѱ��ؙ���!���rS���ͯ���X��d4��+++�Cc]�R0�^LJq�C��ժ���Jʋ�;����F��Ս�s�E�Ԡ��oݵ��܊��T��}("Q�`A ,d<?�o�OޤUt\�6�S�Ϛ��9D\~��ɩ�����c253���27�ˉ�5VTT��3	���ym�������.�l��Ëvu��/%v��@%�98���[,�H9���5!�#�'�l++1�����`�=��-"[+V���J�d�5��JCC��������Cҟl�=!
��������������"�D��A�e���pT�jGF��"P�!d
�@E���6݌���>��������L��zVvs�η��?�=�oM멿�|��ԯ<i�������b`�t���M�͍���uq����O�:���SRx��ׯ�> ��^�f�2�A 7��,<vv_:�{��B��fd|
���ۿ��~NAE�7�£rP �%y�( =������k����޿G���E��s��B��$�����߯�Y[�!,o��ׯ(�1��t�8555�~�
'�	z�����gl�gϓ���h=~vH�&��ڠ�O ��x�2��ϧ�tC5�8��~}����ؗ�P__O�J�j����P'��>[��-,��bH����@�_eNJA�[�!����d X��;
��;���j�L_nRt��]�!�ܟ-k��B��{/��nl��A��
�)ꅑ? U���r� ���Z4��|���^nl�	Iik��\;�v�Ta�.%��M���EQ�zKR�Gx���w���Z�ݽ�7�?G���������e�b�AƢ��a��D.'m���tvv%��F����W�������ހe���IomB�x���[����bT��K��X�ͤ����45J�b���^?(2�7�����W����C!���Zp��#�y0�E����B��&';�%Z=�K�qJ"�`����)@�Y�[�^p6�: k�HH��p�p(��Q��|�<�v�p��x@�n ��@~�u�ݦ��VU��*+L����������#~�/�!�����X����^��f�o����Y/4���������Bhd�a\[� 䚹#��	��լ��^'˓���~�(B���d�����DH@Jd�\g����VlV\��.'˼�}[�6;LKK��<����7��( n�	noN������ٔƧ�GML� l��$˨����\�Cr��o����!·�����#���%��{Q<����v�c���Gm
t�uX�TR^,bd$u�6�/%�\���ɹ��c����9/��� ЏY;9���^W7�O�6p6��dO�ٔ�0�$�fAXS3d�Z���s$|�4��خ�ax������T����mQʮi?z��~��7r�����M78�s�O���I�z���A$Isc��±���r7��:��ؾU�<NY��P�_h����3�@��jż;�9p���1����Zg����=L����B-Ǻ���u�d_F�߆8���� �T�f>�$G��g��fAŹ�����@�B6���޽�ơ�7��nB�v{a8G<쌋��w�'�1�o*`mMNk����nR��mniIFCW���9`l|��E�5�T�'��\�i�a����mj薌2����H�Q���cf@���N㰚�]k�?>^���wp��چ�>@!����Uꙸ��o��%�/j�Y-f�@�7�4��j��Cj*�`.�'II}�Yobo�N��fn�����Rv��ޭ,��A@ן<�}�{������rMb�y���E���,�0ǉ��I3��ݬ%$q��E{���&8��	@B�h��LB,&#��h�ݱ�a[~��˅�TXx�YO���Ɉq�{���H�q�`�^�B�AX����K��[^J9T"��}�B;~�
t���k�1Th^��lRF�����Ez�.)�Q��AB��MC�h��+��|Y 9!���p��\�F'iy�(�����ݍ>���ޢ�R;�M�:����0`AXtn	��Sg�!��f>X�nJj��PY�^��ٲ�i�(��� z���c�VP�y�C��Oo���y��?��}Y����v�eҺ��]��Q �%#�O/����1�>~~�~�����3J�]WV��d�3M����VnnB�Ģ'��]��i�X>��뀠 hHw��'�R�@����_�I��|�or�)-�344��G�	lj�MC�>\;m�4]CSs�ހ������xp�Tn����0)99/���d��o?o_�w�)E��[-�^� 𣅅ɀ5Z5���V�x2���%%���]�m��女���@_�ô�tU��1��,������&Gn���ps���F�u�+++����a��/�ڊI��.}��=�#�������������ȃR��3�BX'bb���S���\S�q��������ߊ���YY���}�k2}�p�6K�����g/��KH��j������؃y�?�fh���Mx�9��"���V�:T�mB?���n����˗'!!!�U��\˂�&6&/��=	}ڑ���ks�rN�<6ν�..���)�bc����K'Zb�w{fG�:"�\�7m�4��7���onm��_Y������y�wpp�P�����ގ��I�ڡ���Ғ��;�$5uf���򶸢L\צdd���UT��m�@j�GYSk�p���@�/���[v(\����:::{}����	NNNX8�4��r��urޤ�M���5�g�\A\���M�����olj����S����|����g>�~\�����������M�?/�����K�!=���J&`Nzw��Dq/���pM�	�NW%ump����}����ֵ������k)!1���'���=�2rK�g���2�R�"n�0hff�����k�󕯤-$C��998�씭ht�o6{��}�O�AB�����k��"w=]L2���oҸL{o���T^���t�B����R���TP��]�!��@�dWOG�{tV3���?T
"�Nve���K\�e�ߵ�-w��[TU�K'<8�'+*�~���ᶅ�����H�%�:����O��a��|�dH�>�rkQ����<��e�5M��筻��׍1�U��h}r7����ZN��!5044$䌨]���8nE��7����4��P������^^�CW����_�'ff����[>�LuC@Ǫ����oJ~N�%�(~��<��O��[M]]O�IOR�"�Q�~M�Z���Fu]��u&c�5��6��C:MWw��-��Yox`���ȵ:��MP�Y������_ �'���ƭaKK��#��ׯ�.�Ay�O��~�k�e������.\���4d�`y�D��������洀?�7pr�f��*�H��5�6�*�Rd����d�n�b��z�>�'
�i��%�gZծ�7NN����vv�A�JZ:��t8���7�s+]��U�Ύ%0Ud1l\|���U���֔��Û�H�-n/<<�ڳb���ty��o)#AO�{���[���ꫠ����L��|U���: ��/�`~��ˢ�:�C�Z.	y�ϲg���$�O��(�>���I���tr��{�d��j��4x*wkOO����w�Z�Hb����[�E���è�  ݝ�ݡ��t�4,��*�R� �%�%��Jww�K��>�﹞?���Ù�����=sn�3U dRY�H=S������J���o����{�xH����h�����u�Sq�0����\?�d������%34���_,' ��ei0)))���4�ٱ����S��a�-��h�2��99q��~8��L������YN%"TD/���O'k2���l@9����ӈ������c>��
|x��ks�]b�1}�B�F� T��)���6����MW
p*���E{;I�˒)3�tC�� Q�.�� g>qjoi�[�QS_�������9�@�h�(6.iT��mS 9��]wώV�ѭ�=����'Mm�͸�@pnP�֊����U^�����Y�Y#�ǧ��	��[?:����"�~�Ʃ��d���Pu�1��&�}��X������y���Ay&�}�?3�zl���*:����а�-.���~�6�`��~�
lfaI\�p�V4��iGF�����W��0KI�MLJo0wF�3=	�B��{Ft��66hf]��@��=ȥ�vvv5��q���=���CW4 �/�d%�� )����_�������A��怽K�0�����U�FJ��Hs���梩�@�d+ς��I�\	М� ����f�� �~������~�1�)P�Zm�8��j7b�[����h� r�ѯ�w+z`c[��9�����c��F�[f&Z��J*�|�#��_���"����b�_B�n�,���5y�#b,���yR�� O�XU���Uc��V��p&LN�kc��zT�����-�}>9��D�p,��0���viN���
�2 c�=��o�o��f�V�???�ygP�	�d����zq����y׮ˏ�������� ipFZ���'t.�nD'�!�U1"�����J}���u41O��4@�c�cCҒ~m�|��^�gҵ���߳I���z `������<�c����u�%<_�66�����g���7�v�}��5S�o��Pu��>-v\�&x QY,�2�W��>�`�ޅi["�]D$$���/<����ۯ�[�o[II�Ք����V��$� 23�R$5��(��a���ܕW��\�G�ĜOs�]$2/� ?	&�E �m�୰Y�Q�R��JuUU��A+_�������1_��@��+�������oG���,yXQ`>`	Fp��+Q�J�^>[��˫In�-���t'sߊ�#	�l�7���+Z8����2=N��m�Ł�9ڨ�[�����!�T�7��`��h��B��fY�cnI���.סQ��qeii�3�j�ᥓE��Pc3��K[���n�[O��7>5g�X�|x
���x���5i�(}K��O�2l����a��c��Ӓв�f#
�LL�~����O�f�,�hb�^�&���'V��Z����=ɦ�+���F���O�˽qf�UO��5G��ەv�Ťљ�Y�=��'����k��2Pmһ��BY����?�knN�d~k�x��s�O&���/`���1������E'm�
�V��X��ӭy������ד/��{B�J�K���߽~�텋g�Y�<�7��ן��PQQ���E�a�s#R�?�0cF�I��I��cccsȾ��A�+����
���; Z�6��T��˧b�V�s��J���Q��^�(�5��8�++�$}씼B��' ���!�כ���-���>�^ns/�K�')(,|����r�
����gS���[?8���2�UVN����c�wTx!f���"�߭q��i}�}Ğ��Ȁ����}Z���$�ԤC�Pq
�4
Һ�O��'����i��#�������;&VV��D�u\��Po�R���nZ/����-9�#�sD�ĄZ�����$1���#MfV��S `G���~4cψ�3���;9���%� ::!;ӥp���oy�����eP̎��[�?�xO��߷��TQHx��,�ɨ�7F0��g�~�B�zPC�'䇇<�q��l\ �����ݐLL�m����s�a&u�gXg����[G>���Fӭ�x�玣}��Λ�u���i!���k�����dce��2�:I�(|�1<�6�_��hyL�Ƞ�G�A�P_8�����������u���$"Nӵ���J���!0��yq` ���_��r��E�/X�֕�zc0hhh���C2��곍 �QS�VWv�u��il4��~�ɨ��rly)f�� �7{#p
���0O[�4NS�}��2����H����ƵOBjj�߮�����b'i�9�tJ6Mju���?�襏XS!cH��0�ǒ��toho%�UH(����4�����C5
Ī��h�#�����ߢl�B�y<1R5̞���������ell���1�1<bnn�xbk��i=�;�'33�3��+��o�i��0*'P��|,�РE�>�~�eyH�$�^�=;o_`�5:�Au\~7g�U�<憭DDDT���K�Z16��]	Y�W������T��\ d~��6?�ti���H��ga� �:Y�U���JՄk?m���s��1�)?&�l���8�?�\���%�K:FR�`Vd$�z�bOz�-�^�`��9*�W��Niq��* �#�#�	ޏ)mmg71$�@ ����Q�Aq�4�h��ڣ��+#
KL�eP�WOK����҆
�	4d;TSWWWH|�����ɝ�v�����b!ѯ�����m���;��vF�h�������ɝ|�*��-�WBC?�m��VA��ވ����4%%%�������<<�b �!�ݵ�Y#�a<A@M ��	�IDtܐ�Y;�lQ�R��&L/��!H��M�df �GgJxV��b�	h�ExCD�CP3FC��)R�z	ǜ�m.���:���|��ab^�� Ep��G�Wf�^�,r*�R,�O�̽P�oS�b122&gA�!x)_��םor���߅:)�u��z��(�Z�)o2E����	D𒐐09�T�����-Q���ۖ~�$ʄD�����߶�]A(fS%�D�.�����Y@�ayby��ƻ�!"#o<<�tL&-��q�mZ�Xs�UM������g2@(�Ԩ���-���^�С$��q�z;7) ���}7�>45�a��^1fp:�|���vF��8���ٛ��Ԓ�w��	�֮7xMing]H�|��qr�h�59�ܬ�g7�ލ�(
KG������ո.˙�>��VU�/�;c�dkF6y�<g&���i���E뭝��xl�|���j2��y /XM��F������Lf?��h���Z�u��C�����iŗ�W�?���U�J���HN��qpe%�߯Z ϴ;3�B�FU�v �T��aT@�B/�إ2��{ʸ�Fd2����'�p�5���lVTTL�$��}�ԫ��ϯ:*���W9?�����&�$�jx�ʺ�_y3�UXz�g���|�1x����~�ޅ�tk?�*~N�{�X��1I�R����O�@�#nɬp����0lJ�y[M���T����>�����A �k�]�Fl�	����ѓ��������zj12�����Y� ���Z�}����ٱa���_���A'��y�Z����m�00:&֥קrޥ>��6Ϫ����6��.��+��/�
�Ɵ㷟f;�+*�G#�ڬ#��)?���	
��OQ̎��py�4g󌔞�NT���8;hǟ���1a1<%�>��DV�Um��Ic�@�dW�x���z_i����b��5�������U�����皘����J��DYYYkؙ��a�����N�G��1���*��q�4��A��!�A~�oD���A9-��,�V'��<��%����0���F-����y��_�j�psS���s���N(�����wsvrc� �AF1�ů
&�- �p�?�R��+.֋��ZX 8Ʀuumm�k�]a-��87��ނ�Y�����H�{g[�ty�'�8�7�aM_�~{[�#���@z�
3��s�b4Y#E�ߵh	5��tw����1��Q3o����C���7��E_U&xs=^�rZ����!Z�cz�fǲTw^8��T:��4����:o�M�Pbq���XX�ƒK���fx�a�4@����_\;6���+��HӖ���_py�}����Z�	� s�A��|���VͅπR_[/]�e�}S8��⭥�63ӑ�vLN�i{���ӳ.�Z���!S�@2��e�dl�+�ܞ-�{Վ���:e��BC�����GP�m�A�����mER�0p������k $QR2�qF��|h+���p�4�9�w�2?�3
͉σ���z܊���R�^�=2��j!�Fn�R��}���F��]Ԟ��j�83���`��4�����_�Tkiy��ܽ /�@ۅ(�69w?'� e�o$-�`xh���%`�'|����?��[X]�������mij�bb��=GDBf٨����q6+Mh�xx�협D�uO$��h��p��^�OkN�D�1�(_�:���,��;��}q=GsK�'��?1��I���&+���.�Qh��x/e
��U��e>2i6���T���ۢ��8Y\.���u.7�Z���Q�JAAA�_�D��{��&}C8���{S:`J
�3�J�Y��"�� yy�ɎS�O#���~�
mې0 �*W��|dg,�/�Cl8�] ���h��
�0�V������A�]�J'�?�����!���[�Ε��?���䌖�m-����u���Ù�����=�����*̈́���C69'��c��Z�x9O��#��R�D��N�3�Ǳ,�s�C�?��v�����@�·���||l
�KPc�}aG�B�j�~��恏WU�F��y�>�WV�‱�y~|��ް.�c�>SA%0�n�P�&i9���N��"�0x1�c�֎���9����NxS쓷ƑG�C��nc�[ÿ��f�NJa:���Sܜ��'xb]�6! /�&���Ma��S��ݺ�� �\��0� �1v�DK�ۜ�����]f�p������U�;��,r���u,~2;�Y���I9��ccJG�vq�8�
۷�����*�Y����]x��Y�O���%�0@D�Ku7GW�����Q�\b�N�52E������VҜ�'��=M���X�� vhS<�S�fd7�}�X�	ɼl�u.�q"Q~	J�E�0�����eMCG��MzL[��[
�����KA߂������d9j�]]'�<�|��'��C���+g`7��F���xf�����G�k�ߴ��%T�zjk��_��0L][�/�zEFERl��Wͼ~�uM\~�����.�Nw�[�����e������V�����ھ^>%��ż=��qT��_�m`��V-�װ} �<W�O�L�dc����7]��.�:����[~⠅���:��� ��x��,���ot�y4_G�z6�����C��gL���"��*pm %筈��3�ۘ���j��}���3'�$-�/����'Bi�d���'慦���
~��^[�zJ.fgZ�������Nj�������l �U��MY&��2�������c�)�i_~�������H>U���V�ue$�����P}x��&89�����=*�F�f��g2{}C�X\b��fu�u��UI�~�I�;��]�G'th�Ͼ���B��j�5�v
i��G}�c�"���#����@#D�����ݎ�O��ݒ!f6�چ}L��:zz_�3��s_�"~~�4
��G��4���j�C��R?��}���쯕N_�1�[�Q ;dcdD�"d�~�j�JT^խ�t����իW�Y���z��-�`����©�4Q��q�j}q���:������-�m�gM-��_��^I�җ�A�+1�9)�.;��OH��4�f��g�q�XM����~546n�
����UTVv�JAf�c+Jv��ܝ	��W�ܸ�JGG1��������|������[���1q%�g,�N�N9�'d-���A�m���nN��<<8��������U7��st�$�#�çܻ�蜦����E��^1����_���`4�~�����p�)baa)d��><�l��/B�)��������N�̜�qWW��@�n�S��3%h$uܲ��l�K�����>W��{h�5���AE��%�����r� �#��i��i���۠:l�G@ ��,�,q|��HN�vo;nO?��I��Y��� �T�ϻ?VNVZ�66X�=��҂�:�.��1������xn1o:s���D��8d��r�>���?�P ��͖U��w"��Eq%V��c7��a�B9 �q�IcɄ&&U�6d|\�v�ˏ@�f<�4bl������B��~27�Ce��~���[Ef2q��b��@�f�>=\l�+�@,sJ�Wz���ޞ]^tGh |�c>f;={U���r���?A/�G����X_o)z����1���z�G=�	����̗�������?���^r|Q��y��{�!(��Ůf�F��隐�����2AE;���5ZkH��Xj3���k�D�\}����,č����x����qr�|�l��1;�r�ĉ��7�����/�d��d���4G�O��[�n�c6՛M��K��T-�F��L��FKR,�������MM $�H�u,��ؼ�q=c4)V���\N
qE]����~"� ����1����{8���W��n�b�k0ך�ZƎ�E����v~���B\%��,�^r;��@B�d�ޥC+�.ʏxx�q���Z���B���=49[-T�N�/����x�����t�ƶyz{ݜ��E���Xli�}�h�ҝ.�ll@^�k�"!i��:�p���6���v��"���6f�G>������R�Y'���&��:s���<��ӄ��YJR��ĖB[�m�Ll�e��~�̿�_�Og�
p�<x��L%'��\�����VnLM]��l.L�?QӰ�7
\_j�+1Z%�ǧ�OMO3y>���<ٝ��t>�aK��g����HorJ�;���v���/H�`3k�~}�Bۛ���t�[���H���:�ퟚ��s7"����Ld�!��H�k3���+R�1�ax��.S�Ү>���i��>>5����]�S(���T[[+�ˠ��@U��(($�l��!�+�B�E����I�cl��7cׁ�Oa�0@��%���I��I�842�;�Z��fꏮ����2R��43n�7���s}g蘬��3����偷H�a��Yh�o�5*��6;\n�؍Zz�Ņ�d��#3�d���пR����%��ϲg��d�BV����S��4x�g�˵�Øz�	GFF�-.��TC;$7��v<5�!���C�}V��x�����F�hz�^������W�h��{)ă�r�I��߿/2��͒�5>�Œ�����i+*�L������(c\X �g;��׹b{����J0�9c�T[V�����P�o�5�v;�b��DiWy�<կ�є���j���`��bHJ@9�]�Yj�4���)�A�/�˞�|�����Z�����f�1dL䟆������1���[�Rwk�̑VǲT˵ؔ�W�Hvc�\�[q��D<��/,�-K�E�3��|a�,Oj��~��hQ�_Z=0V�����²�9[3�	f;{�q<��������I��!ss�$�����iks�[[[^@'��WF��ģ~��8�PS			H���Y]�:CSN�xy]�)��o:�����ZF��^��Ȉ���}9ܚ�>X� �j�f�ѕ��_V�d�'����˞��s����q� nA���xI��D�iV��j�����q4��P������;&�T/�Y�!f)��G�2�
FQߢ:��}wXd?;�Z�l/��<<�+��]ʇHm�Bw��˝��:O���K;�!c��o�cߑW0�t{�_O+;o�h*�����V��/ug�����w�e���o��f��4&f�&c�a�\�z����x��$(�u��mT�(�y����v+�����.�O&��|�X�	c�㶻qک�6�ދUI�}�֩���~��[�0s��L��$�t��<���:~(s�geaA�E�N�����3�6/?��,�����]�㢖 ���`o�ŲfA���kf&Y�fI?���޿��i��������>8�Dfgg�g��ɢ5/�f���P���>��I��*{m��IVk��=��Ӌ��F��H�t������8���Ɗ��Wo��7���[=�r>2�p�.��E�z������פ����[(wg��YzA%!A�]�8Ve����Fw7BL�p;�e��ap��-����d^��.��Ϣ	������M�^�	��1B���~�/<�&�������R�P�4�4 p�D�b�1�s��*�8¨���¨�Sj�w""���K��Q��a�ynZ�i�����F=�O]5�߇w�p��E8�3{w?85��AL��ʖ����7�����a�.��}ao�r�8
��ĵ��ӌYG�����A��'�Dt��su7�^�7i�������Q��q���a�Y�]�����o0>��y��nX��wy4�h�n8�'���̼4�YQp��8JU*���K��jy��ϟ?��︭6�[u�l�X?
�.�&n���T�\F�������C������1#����)TI���W��N*MoR���wed	�b>���Լ(2(����2q���4�!3�V{;C�:�C�v����L�Yi6�OZ(��wD[BN�gm<���&#��e����5�yvs��=L4��FG����()b�%*��'D䨕�=�]͖	����ei����0)�xX��}.�<M�h�m�+)Ezΰ�LI������Z���-V͵��Q�3�8�A!JĨ�9��"�T�d`�Go��:����/��a�%�#Js�����C�;ˮa�ۉ)�&
�������OV����0�׵��}i��NŽ}֘�y��$*���w��c�ii��<wP�H�n�^��=ۣi�Ȭ
���4ٹ����ѷ�4[?S옕)�g�U	����Lj��s��g	�x� P�YS��N���9;�~�C;Vb��}�nHh4}o)$��
>>��h漶����]H���k�+��FA�?�T�:��om����=%�&���Fi��EEE{�Έ�`�t`�w8PM��z"��8��r
��c),T3�ҸP6�+?���ɢφ=W8��\U5Y��{�M�Ǣ2�*�p7O��a��<h�m��^(n����b��KJ�4<���v�h=�QJ�N��
��O�F#H�g�G峮)�^�"����$�;��S8���IFX�Rsr�:+y��=VVtZ�]Zzv3j<F���_���]Lsَ���� ��j�[��m����G�dȌ��������s,��f���Q��~�+�y�_�2
͊cG�)(e�$��u�Ʋ���ķ���B��Q�;����j۶�/�~;?"� |+� ���z���������'�YrX.�,ax����WR��i-����v�.I(KJ5*~�r��3�]�p���UaJ��.�u�f�A!���縜WFF�^iM0'�ć��}��s�_��v��;2��x�2��U�А�Bbb4V�ϡw	~���1���ջ�����C�� {��y��� �G}�#}�����������k�Y:/�ϔ T\FGF���B�@K�{�a��W��J̝dP����ժ��������$��5�����w�'��PWux�wC*%Nw�SM���h�����9M�>����A����ʦO�?G��^�%��Kj�hJ�ã��&p;���\{ �UZBv�c9q �%�AYMpo�ؑrND�i
��Z@	����Іa�8��ۏ��3~0{W�����ޞ���eF�=ߏ��)����5ɞ2�T~it$=���	��4������a���h#U,��*��{��/ez0���>�e�SE�dy[�9E����<���?w��:少���/������D 0%�+w�����p\�AGG�=it1'T���0(xxxTiv�h���M4GE�x�onm5��'�����˱~���f��):?��8���S�Ⱥx�0-�+��n��;�n��IDH��q�Ǭ�����崀��v;Y&s�D )dEr���vt�I���ֻ��{��'������c��, �t�hۗ��p�����:	d�s$��{ͥ����zz$�9Ġ��$jj"+�A[I�Y�n;r"�B/|&f0�aL�qOD:S����5^h���[�U	��v��=�E.ͭ�]h�o��p�h����%jN�o��R =M.:�sIܻ��t�8����U#)�%_�\�H��m���pʍ�-Z�ݡ�Υ5HM��Ӑ�t���	�#"��W]��d�gkBAE��N��e�/,v�1^��ü�_D�a���ߌ����M TB��H���xx>v>i���|Tow��|��aR:����t)��ƥ��H����k}<<<+�2944�GH��SM����Y@�b�Ｉ� �l�I;���i�-<�'T�k���<"�@�j8J���}A4�%  ������t��;��~�:%[/g? ��;v��]�y? vV�8I=�����q]/w˭:`"��7$�����F���|%%�J����F�63�?00�o�611�U�s�g�v	qq�����f�X���b!���Q�c��ҹ�a���|L���FG�c�=Y�%wZ�W��wQ�S� d^<��3�qp`�7���w�%ܿ��i+
xEī|�Ⴃ�������Ԡ��C॔J�['!!�_Sɷ�f�_���+��l��*.�����E06���p2���p}X=�q0]nv�)D������
��j����U�Ez��"|no�3k�̹+tj�����Dp�����v;�����E�������u[u{�����Gy��(����>a ��� ��{w����!��M�x�a�5����j��
~#V���fE>��T����Iؘ��7F9<����j�q�\@'�~n���`����R�ن�,>3s$ڈG�S�Kr��\{�J��;JJ����?�I�(va��2��ن�q�|�Ng�\��W�Z0�7�4��� �N素�����Єc?mg�i�������Nj�+� qxu���

+���V��}���{�Xݹ1�/�RFS��	�k|��R&�������W&���x�Ϧ������]nP몛-]�PtW��UT6G��(]
��}��b��t���# =�!��/�	^�����*Jkk>]�1�'gdDʧp��D�&��}u],�ևI)�����]���ugb"�m^^^��8M�����@b ސ7?����j�}�E�^Q�~�v���PLu�o�L�j�����,-�,�xj|�t����+=�0����X��$x���=�o�戻kL̽�A/h��H�l�{��G:��S		L7���`�ؽ���1����F���� ź~h�9v=��C'�qvD\l�����Vә�b��I�Jg�?h�6_ƛQ*����T��Qڡ�6P���=�/�߽L��ݝ7E��7pE�:v>)��|]�� �/Ǟbf��*��)QQQ�[r��cX���V�n��>Fs�,�?
�B䴜p&��#⤤�#i�Uoӝ<<BSR���B$U���?>_-�W)��u��~�N�433C�%\@j��jm��};�V��{q�Q���ڞ�z�@����M��.�h�6��
�h���XVP\�r�@A�Ì�l ������+6��i�Wq/	8�Vp5RL���j˥Ye�{{g�Fԏ2�rl��J9�n���GPȏg��,���vw�Yܧ�𽺀��وh���,��qM�J����E��X@AA'I�ڞGN��q�vG�/��O��FFxߛ������a�A�|n�f�t�si&C���2W2zoL`�<��Z�ĞB����]R��������C�ۏ�\ ]F2$���ED�H��.-���dw50�)�}C9�.qxQ}�|��E�Y� ���c��v��{<��?�bg�4�܃T�c����J��98T�9�fO�.6�lll8q^�zA�n���yv
�g�Qȿ�{eV'K���!fm���
;��R{�����5`��p=N+o�[�����h"�			J�������e�o�Ym����.Q�ʠ5�F���"�#'q�[�/��� ��Ǟ��c�>��*�J��Q�ZJ�R�Q�#��[��0iV����ىrz???N��_�L�oaX{��?Ž_�E����d�����(�����������ⶏ���_~~/`?����,KGO�h;[����������3l�1�������xC1��|Q�p��\��]��QaPKZQ�uK{x��d׍��+�>���7�B�]�N�Ji�V���߬�H��V�Z��م��LL�}��>���.���EDD�c��F�L�J��U�u �n��(k����ZZZ��ܔН1��s#q �LLLREً989��L�.�i[q��Y�^|F�"�Ѝ(�s��uB
n��ƾ��;��fd�Xq�B;�� 8���G��oA��O��M.���f%���z������'��>�����'m�p�����h��d�jLH�v��6�2��~�@�	�L���[�=�a���Ó�X�B�*@8��n������@�~/U��p9t���<�58Ik��p۟)�_�� #�~�����RVR eR�?<x�o�a��
	��w��o��Yj%�U]:��s{��	����XGω�g�.~�"����a�Jo���,�q�T�����5�{��x��^<�b��EDD���Z�������v(��`��8 .km};�E��+�R9I��x^�&�$
�c���Tkb��s IQ�;iij�����D�4�^ZZ4XR��L��0���W�a��"�娤��~{���� �z�b�t���Xc}##��u�.�g��הkgP��^��"��Oڎ)��8#E�����{܈I}�ݬ��h.^=>��E������b,@ɶ�E1L��[�K������Uu�x�ؼ^%#�c �B������q^�01�1A�@���­8��� ��#^�@C�7���E�RG�������4�Ǎ>t2a���x�p��_��B|�^��/�Ȍ��vq�.n��.��l�|AC���n뤁K6������Y#�Ju�/L	������BFmm���6|*�fH4�9x� ��t2��Hv�DO�ty�?�e��f�4���3��99kO��>W��Ty������`�!���^� x�2\y�Ls|%LDB_Gg�5�ڻ����nwl�\�M�T�5���A�!P�`)��|L��V�}5f�^Jq�p}Gg��J]���D�4-=�t��7'OO�kFz4�����TU�3˅Tzz�s���rrh4ק��R�##��f�Tqr?��~��R�"e0���\�23���l��i\k�#,T͎Ȋ@�{��l��a�xg�����i�)��-�[��m��S�����i>|aH��[y?�3W���;��xz������f�΅�[qQ5���x竑���,�K�8X�q�-+/ov������-M,���=f�X_���^�&�~��)�}ɋg
�XY�Վ��Mp����N�8|%#WD2���p��N��e�c�8}�#S�1铭��� 6��w]IX�/KF@@�iIz��bS�z��HLNIdT�eYmHא-n��I
�==��}��7�_�0��V�rU���'��^���CjZ����4sM{�������xR��h�47��mhW�o�bFH�xy{�~���2��g�1�%|����ES^��s} Hҳ�@R)��i�·�K�3����R����!��R0@��Ԕo:� �rejji&f�Y��ڂ��Y)G��Ԭ�����3�3m=�@�5���u��]&���Ƥ��/姕��r�,b�@!L���󽒜)�����	��@E���Qt���7O�qq�� r�D��ŷ� hA��5�voj7��\V����_- ���j%�?a���v��
]b.��8�����e����P��{V�����ݱ�'tx��c��(3�K_e�(��r�Vl{G����)����{��sE�)%EEK�2!�ߌ��3��=�4�o8�x����\m�B��k�Z�ќ������b�ˋ;T��D�:�����*e	F �������J[�����y�1������6�$���|����ؙ�^V��b����AB�տ��֞^}�s��"$�����c��j(��
0\ݓ�����2�K���`/�1��J�:1ɾ�P*����$j|g>���
?ۣ`ʌ���ڿG�@s-�K������ Ƙ��a��;w<<<'dA2�in)�D}Z�f�܉`{z��#�k;^WǢI/ G��C��c(CJ�ʶˀ*)����<nb���!�k�u|/8����<5r��Af7hc2�8���s4Q�_�~��g�7����}�R5z��=��uF��0|�7o��#�g+{<W!"��I���Pc܅����,-����5*��u�Q�I��'a֪(��҉s܋t�����و�������gI*��~Xnq?��W�A,��<]�f`@�/�(UC�\>����|����S�\I$�B�mG���:��@�~x��*�^�۽E�TwkSĕ�� ��� �lv��w�i_0������tl/6�� �RbFݼ�-A�0U�S�ަ�>}k˜��� ����S0�pL6�>�����oΖ������8��i:33��)X���n�{k{{��c8`����, �#~��.����
N�nyd��A^k��q������<�H�e6�0��O�4�Jp�g)5S22r�?�.��Ў��Mako������sD�g�Q��r7+:��q��d�$�L�<����p�'H:�>`�z�;h�F|j�Wrr��W٩�?�Α.��]__��u�Y�]@���,J�-X��F�e�5g�՗�K���Y{��,ZR�E�n$��^�8=��0�u|Nd|�@�����x�o��^�Z�(;�|�)V>|$+�����E��&淛Dҁ�ҎRv�~*��������Rs�cG�[����
|=O���x��IUut���{��@��s2��GG��<�{b��y���{�7�#^�/���rL.�|%�,���,��0?��̈+{���\Q�����c��Z+�	�#Ɏ/�x�����Ft�I�H�񍾚�Z.7��7��	������0�:���P5d�+t�f��!��3�Z��y�:�ߍ�d���r\���>^�h�V�HM�ny⻋��D�y-l�%��+[��0���>+�wi�i��B�-����,�S�=��uji�����Ly���11���7��]�HP(Zh�%�����q����v��-d���
��_j�r>�D���ds�K�]�5�>� )Liׁ��4Ow��>��D�©:Wi���V�}}$���K�uX	���+�K^���u���H4l�>��V-s��!|���J.���d��9�7�sB��$0�6�\g�=�ߞ��' ~��7�˘�<&�qЫ�#�`+�zR��V���2���s����=--�j���>�e}�r�x��vL�vt4r�^7nYKe����1:Nwƀ�~�
ͥJ�T��e�}*�"Wq��	v�	����f��M�Z� � �Հ97H�ň�0o��v�mmҼv�����0`��t8�˙�u� �-4��[ZZ��Ձ�<����VN���A�ú>̫�cbpꆿB%�%0��O�)i�p��j����㠽^��"M<g�Q�O6���#���RW�cǸi�	��os��/�E�x[�[�T?ܚ���ip#65kQ�cN�s�}Ī �z�YeP�&I?�\Z:h�mDHw��]Yɞ������|����E��	P?\��nAo6��J@��=���6�+v)dl,v^)�(T�Y/TNk��)k�6wi��L.|Ua�(i��{�� ���
�XWA��~ZU�C_���	�A�>��9a�k.P{����C���Sr�k���V����n� ��Ӯ��NK-o�-�Q[T!ƏI�R6�:�h/eQǥ>jk��Jk��_�P��n�{�^o=���ڊN@�P��x�L������\9�M6�ə�B������1� ]��o���).[1VV��{udd�EL�4�*^P�u՚�3D�N_���n�'�r��]��cvo�0�ݘ��:݈��ϧK����w�c��W)�0Y��d�N ���QRk�Ze�$��f�w�Q���A�ջ�_#�ٹܘǿB0��X�"�# �s�|�k�pX�1�J�'!1a�ę����̰]�Y�j䈔Ӊ��_��A���\B�D��z�禽��	/�$˗�-�d�����|VT��p䍕Ѣ���A pW�d���z
	e9k9�,(���O���v�|r������_Bǯ!�0O ��S;Db �b��$n�S@���w:�D"�ݳ ��w��� 1��b����"0���^_��@������>	�6{"5����pq��+ܢ1��9��{Xp1N"�0�h����#ʛ�?��^ ����������^�4z\ʇW���+8�Z��Z�O./6�tz?��K2峷�r�@���d�:�l�8ɋ���Չ�����Ș���������@n��Sx���?�zG!6�L����c�i3s�61��[-b
u��{z{�b�� �M,�̦����?:�1��9�<�hhl��6>���R����)�v���L�u�xw?��̊��{��&���C�S��]	c�E��6q�]]]�Pʹ_jj��\����5�/��~_�l���,���Z�lº����� Ǒ����	�e-�4����W[M�?J]��(�B)nŽ��Vܡ��K�Fqh�x�R�-H�P�hpA����~��{�u���u��5$�g��#3���M,/é�K�9�f��u/J�0��Rj�8�?1�K�֣����òӄ�Dn/�\Sn+����HɗD�k��-럹)��y�՟jbb�A���[w��<E�+&�%ց�Y-\:`�k�W�y�z�l����PqoG��sy�3��Mϩ�D?�p�&Oc��ϟW���*V���&�z#������S0oS�2rP[��[r�zz�dnbw����e�GB^�Ł�%pޛ���1��,��-buX-_|@��>`�ٸ_�9r��d�odll����	�a��������޾I9�g{�_SSٜy��P�Zi򺌼FDtUF�"�Z4�	d��}��$�'��4s��.G��˭�z+�=��hJnOVSSǧ�Lr_up#�S�ی�=�H������@�\l5�/�~�:���[�yU&Ӹ�v��h�R̠�@��#){pc�;�Hd*짴u~~~���թ3(ǠQ�4>�IN�n���<�cc$T��e��c��mL��v�����Dt2�LL��]�j�����D���39����#�Gs$�/��!+����N$l���#�H9��(Z�
w�>��+Д�$�v���b���O�Z��R�_���"K<��Y\0��"��[~��9وhm�*��6D�vGQ7��Q���ׁ:>6�Ҙ��u2v>���G��y^�w�}�c&,y�dn:co%]���]y�ZV������2��Q�DQ+>jq�,U��K���C���*|͂�E�F��:V{���#���$�s��q��҃i���*�.��
�v�0b9Kx�tۭp��Y\��kِfS5mi�@��Y� ����mm��$��@��ᩐ?���Jo������V\�Bcb+_ )�E��.�occC��x�9�:Tu/W4�X<Sљc��N[�Ԉ
pWۜϣ���!O�3����=e`���V�)Ӎt+��+ϸIlF�vښ��]���>]�ݿruޡ�V��9������@����M�504,W��3҇�Z�'��@ z������s�c �;-���!x���6(W��O �A�����Z�Ee�p�
I����= W+�l7S������C��ϖ���x��B9���;D��J��Ik�������%�������'j;����f&�vzA��B�>��f
ʔ[|'S��/�o�EMS ���r�[W?��Z����
ת<7F��uz��e"Rd�L!��PB�a�u��U�b�*�ze��3���!�R�۷rI�`O�d���(W���33k�Q���Z5K�6{v����N�&sO�]���(A�q�Y�ȅ��T�YY�G2k���?KKUP�C[y��>X�Gj*�XɃ$r��Q9���D$������b�*�r�/�"���<96y9��B�!YK��~�zo���c�[p�գa�_�􅼡��r�����,S�X�@�rzhbDJ=��!:��SZ�����"+�yd������YGO����f^�Tx�y�x�آ���� ��˼��u�~Y��\��gٰ� ��+)��o&%Ój+>��2.
���&n�H�D�7�������}} V�D�������ҡ�E%��M��V%��f*��?��i��_$ke�ǁ�VU��M�.�����������f-'c����3����7Q𚧧�͐V�������y���zȯ}�}ހ��`�}�\9U�}�n�׍��I���8�y�ˋ:x��[���b�X�� �8-7t"�S�������f�*�R��7�/��n������T-����p�r�̓W�R��i���s�s���pi�>D�&!>�۞T}鶄;nR��篘sג��NM�� Wv1�~�j���*0��������_�U�<���3'9���7~���� �
��-�J3��<���^z�OD>e}�E����@G�v�C<0Mm�X�����dW������� �?+�ؓ�#�11�����9�2�Ͳ��l�K��!�E�7�j���'��\R@�|���f�������w�q��Ɔ������X�'�~�� �t���l=X����EWO��J��Y�T�b����>�������\~��YQ���|�Y�ʩB@�%�7ޒ����i��ȶ�6P�|���:`�W�@�0��7:���
7]X�MK{�ZG�`�+F�0ƖZW��"�ȗ��ގJ��0Ǚ�����q� �DY��E���\Щ ^���;B�m}�����J?�SZ��^�mm]�/`���ޱ�O�1V�
�+#��r�<��ܜ�!���<>�.����}���9�:YHJKH9`���:QN���)�)((x�07��3�+__!�:kZ�os|%U,HPDT�F�J/�����������p���"�߷=+m�K�~غv[YX��D�S*��&��~;�{���F���2�-��ܟ���V\�\y�tX%������I9�w���P	�_$E����M�f����2��:�u���y���O+��L�nި�L��ӳ�7Q�����N����Sz++{U��Vf�P�����O��=3U�bbi��?[Z$�k�ɴ.ι��7���|�ż/�aS��i�N�a8����ln>��"�,f���|�I�H�2F��,���Ȕ������Qu��5�gcl����9���G\���'n# l���ǳEX�3200@�;mz�n#�l���_�����mjoww�,��=�6�bFp�|��΢�ԣ���*GǨ��3γ����F��'�B�f��踱��~***.ˍ'��_e�d�8)>�_h���"�j<ܝ�Th�0f���n�</�k7�@��~�yp4��;�a��w��n `���9��ΐ�4_��W��:�Hq�5ɢ��?�ו�y��Z9��e-��x�_q�جQHn�7&"�O5��m
�s���f�)z3�=Z�+��UW6��c?�U7���Z�#�(J1����Q���\]˜h�_g�=/�;�^�O�L��B+��o<K��z�I_UV����V�IF�מ��2o�����$,N_�S��t-Ȫ�?�#���W�O�f෍�2Ne�����!mmo�Mǃ��K�f�p�h�Χ�\*?����A_���(�M�g��!���)��av��y�'�އ�޼q����������ba�Xiru��������lȱO�)���Պ�����pB������t�t]�bcc]������,v/�P����?}��[>[-��;y�K���J����ޡC������q k��Ύ���8!to��`�	8
W>�A����K�ջ� yܼ�<�r&�X[�ZYYљ��E��S�?��v����m���8)���X@XW��m���1��#4br�r�n159I��H$��{���jo�Z�=a�Dtu�1VL)tI���$��L�.�I@�7�u�LL��۪�-S&��wֺ	�����-\I�S�(���P�lq�;������v<̣=/ݥO@bnER	����A�y��(#Ϡ����^�m	NnnI'�*g��r�_R��E9n*M�)t���ǔ��B� ��S�2�N�����v��y�]\\|$_]��+����ׯ��v�L�j�&���	��!9���섄+��6�����**�~�_�h����{�	Lx*.���z�W������SP�VVJ���ϸ`�'q�/�cJ�YjLW�N�NK�`����][��.�-7,ӣ�	��,��P�EC(�� vȩ�i����^:���{��UTT�k��&8����9�����ot3�Y�jǞ����\>��d���m�䏎i��Í�x��:�̞�>^
����`�߸cVv��T��Z�A������e(�< ��!�: |�ѝ������fa,��4m���/_
l��c;U6M˟,2D��P�:L�'�����{z`j@K;񈼑��q4.ވm�w{���WX���%�$��V��4n6��j�0QkBWY*IN�m4�����&|kBK��Փ`��+b��:�#�S���n+�����Blw���=|�5#ؼ�Hhoo?��x-��_�ϒk��	����].��H� ���;%F�nR��߽���ř�D���S�Ne-��]��>�eH\��eD�y��c߃���BG���	t�2y�W����V�eấ1H��t+'L|BB0�~5癐��x,W�~w�s�޽i]G����v��~�^8�pK���(�6Z�ٳG_Ě`�<z�������#����?4��珬���]r�g_��҃pһ�V@ُ��k$O����T$|@�zt��+���r��ܪ+pg�%H�&@���	�DBb�9�p��b
�|���ٖ��Lh5�OOM7��L��}t�NI#(y�3����.�����,�ۨ?{
��f�|ߔt��=|�=���hq�~��
��P�"$��ݾ���e�^!1h�0�/��# �-�V�SqKIUѹ*`��=6��'���m��>a�����Hn��A�I�+�r�}L�߸-�F����ㅡl��@N6�i���&ץh�L�m��g�=�G����&��wQ~��d3�~�8��rz���@����5��yhnV�0B�M�HH�l�K����6w�~.o��NuP���n�ȕ$�Yg�ً�����=����;gn��z&�2��^>��+��V���B����}�����֘���rj�u��D�����C�dW�yWEA(�(b$q��Ʃo�7$:�����łO�β?�.o5������6�}C耽�\\\,��^-~i~���K�L��4��25�헖YǞ/��m^1>�B�f
7��B|��xU��3���H�ͩ|H/���X�M���U��MS��ZҚ�p�ٓ	�D��P�X�>S���.��#����s�]�����VW�&mJ�Ǚ+�#���~�%���̂Ov���\m��xw(E%��j�n̞`�O:�q����Z�ș�k�w�}�v����K���@���ɳ ��k��~��J(��5�
��d�%*;�4�ڽ���G�/������e��yp�k:"k�j�%No���HP�Tn}�eZ�q�i���H`�!��4������|��B�	�^K��ݒfSQ�QOB�J��M6���w;JpsD�v/���H��B�}~��NcQJ�[��TV��{a�ܻ��.;�� �;����S�9X�D��T��A���L�~�a����=����X�IH�O�zYY��ߧ�|?Y[P���S浢�b�Mv|�[�3e��&��z�՛S��T��~��SSS�;G�mD,�|�� ���Y�w��jfgĘ����%Y܆^5Ӈ�J��޽u.�负({6�R+��Ғ��[��X����~�,"3B��}�fX��>��A�����o<U>r3
<�,p.L���4��v`�Z̔����*乑��~��졿r�k��꠮G�fq��!l)5�g�~|��MMz�냕 �[mp�6'2ECH�֖���_�! �(���������KK&ꩅ��rr]��b�!�%�%�TM��qeF��?�]�]�v��{^	��)�0 &���y��Ը	��;���D���]�SQ���|w�����B������2 k|���yu ����Hޱ�0teY�{���i��6=������K5|�h���({����c����M�k�M��]vcE;.qD�퉻�V�w��� ���~C����;x<��QMŒ��^͊��Oܑ���~s���R��Z��C�2�'�����{���}�p�����l���3p;���� ϛ&��q���]��y��\5�e�h�v����c1u�͇�᜵�:��n�5�L®(*�\��AQ��E@%v����n��k�!��"߄L�(�w�	����+m����/��b*o��y���e�}5ğ'eg��&���iY����zR��i����ך:]�{yD����E(@��~Sgw�wդ��5/�����ϝ�21m	Է�v�6��J�}��4�����������'��KXH�+���fVM��Sh*j>��1�c�GC���1��ɬ��#c���Z;r�������o x���IH��杓S�,ė��b�Z�X�خ����kx�ٸ��<۴��0�"����+�5g�@q��njiiY��qQz��3�X*�=�$ �z�.$�s�WHh�늻w�z"f*P��o\�(�_:��Pu1���|�c:�6�v�;%Ν��Jd�k�'�FC1s��<l[�������E�V�������g?��W�!�Uz��	�����L�[+*�4n�_���I���{|�ɛR�W��~�?M���;��#"}�� ctTq.SP�l�0�̭`|����;�֬������Ӄ�ś30���be��T^{�޾ ����Ɔ}3IuTX�ܳO|�GhTvj����Tէ�FQ@t�����f�2
R�^���6�to���к��'�iI��y3�3`��1��b��������Jj��&f�g+/���V�[�lo{�5��!)9'΀�WX4����]�Ӱ`%9�Y|����==�������u�r��~���?`�`�c�ЯM\x7J���M�z��Jւ�Z,�^!}4��r�_��f��'�N>-��R���o�o�/�9o$^Ly����nA�����y���{4z�|k�*�9�|U�O�����LY���V�~��/�R���ϟ��a�bK�b?7P��鳥{`��+'��R��gʸ#O����/���g�_X�5و#��1PO�7�֧�eF�-�O1jn��zx�=a�S�N(f8�9==�i/�cF2��z����o?�L�1lڏ�yu|r��2n��/&o�T)z�^��?r+�e0\Ͷ6V\�ܛ��D��
-Fq��c
S^27^-@j'�xzzZO��jU�:������X��{����Hv{eNN�2���X�v!9q}U���c�����V����ҬW�
���y	���\D]�hi���G媤1F�����4�aO7�5�'u�Xր��Bm�����==�!����5W�+���}�AH�/���		��΢X4�\D��&�v�0�nih�����vs�7˼�r�c�1��8���ѷw' (Ŵ�7 c�S�3e�Ƽ$vI�x�2MC;M<����(�"2��}wk9?B�P��sl�!��_��>�zP�<�ՠ���Ӛ�TU8���f��%��s��E����o����z]������l�
��*��&!�
�����K�I2C����P��LP��9�XXu(%�N�Rc���8��b�)�&T��6��܄	��-�cK�D��J�
}#��y��4��N���G~��E� ��� 	\�,�כֿ�2�޿�)�{�$rQUS^��%"-����ͣ4.O�����p�K�6�v��y�͔���M�?���*�G��1�!)$�2W%�e�+3��:wz�6���
�t1�w��9̭6���5),�n�;�+����,��-����c�愻NQ�{"��]�V��66䍈�A�(�i~��%y�����-���`�/e��-�|{�l;�ВҰ_�-S���H�{Wgoi}�59A���Ʈ�~)�I��q́+kwW�B+-YR���m��V^$�r}��H�=�*�!��du�ʇ��HPp�=X���u��vgQ ��$���xHM���U�7Ml��*����no�)�	d�t3���ı�y��]����pg�M)uG��̹wA+*J%��2�$.N�+l8���ֻw|�-p�3�dW��p�)[�f��|�n��DU�aܛt=���RRH�N|>�7�%L��-B��䪻�{˼g�92j�Μ0|�9��gi�p2^^�}F��e��k���������^B>}�	(�r�?��qB�`/�|��7T�]W��>;dSN��ja��`ׇڇ���3�+YZ���m�_�=�Mq������0o��M���F?c~�^2� K�����م�RIQ��<��!<Ec~k����+U�biiy�^��s �Ԩ�8޹U�<��1��=�Aq�_���^_�˾���|�{��
8\K1��1:�����dŃVV����j$�����Tf~����7*����㢒�p��Osa\��BW_���Q�rT���̵pK��q��V�������e|F�E�#?�����#ǔվ��̑�SS�K���2-b��|o��z�W�=b�>{�X���pf�&<Uج����ɧq�F���jV��������j7Q��jý�Fw:�K��:F
�KKP�_,6*�[����"_�]jb�#��1�l����"�$����(�"��hss�G�<��o��O�]���
��ٜh6e�DP�b��[O�V��Q([������˱�cV��7P�������u�7k��g�jy]?��^��ʒ;GI���_��\���J8m7�/,�o3d�lg���E�7Q!m�y#��*`��Ru>z(�ON����UU���Xw_�$�/Ymo�J�����4������Em"+e
[� N�$Uo8�I�7TPPh�ԯ�j�a�z�'a��D�_1��W3�+M�����N]	(0�� �Q'�8R���'M�0����� ��+;aA��G������Q8��kV��^a����ޘ��^J���TJd3���;b��6�"^�. DZ��f�~9	���O__�X��A@ZO;W��`�������S�|�\B���I!س���\���5�!(����\��pI�(K�t^�Gn�en��y�W�i��w�g�޾}_������i�"FGQQ���<�_jP�})���*@�%-_�{�M��D�a_k���u��$�X������C=b��MM�RꯅO�w���[�B���ٍ��:�<٢�E���;G������x�t��)�#ja�.��t��Z�>rz8*���b�#�������ĸ�b$nt҅��k_{�BMD���0AN�/7����̶W����E�p����{.��B�QF%��0xH�i3�b��}��S��~�������d�a�_O��|u���G������O0��΅�v�vC~��ګ�K�ڲ�Էk�j���o� 7:3���F��ќg���W�cF\��0p�N�q��`sZ\��3h��b9���q����4�Y%���6������C3zx�c�:��i���b5dn:�ӊz�/�bkǙ�G�u�G���f�bf��xT��K��w��K�)�)�F�j�b�F���VM���V`��a7��Y&�5�4T�>|}�0�뫇CܱI(ְN/˭T����έ.��$�-ؑ�
e�פ}�G������B�R��F���˄�l��7��� �2��Ӓ�Vy!�ZĢY?�򑑫%�*5�C{睖 |}�
}��/���//�o�]��L�ͷ^�w�ח��nD�U�d�#�>Ym!�i^U�r����%�����h�O�3���.V�p�i,�+l�꿞<h����Z�7�I��ԕ�(s��M_svNTUUMAѫ0�Ȯ3��D90�U*���"?����}�ew#w8g���c�vY��í�c����}��>~#�t�6�^���u>���9�(�Gۿ������=KC�]��0��O7�{��T��P�;�C�{nM�/���Xґn�����$� ����N6K��v�������`��u�R?�E:B _�:w4�P��%�>>������Tl7�W<�8�V�r�j�r��nVi�c�=��j���ؔ��[�$�Nd0�Yhǟ]�A�f�)��x�gӯ���`Q_K�,q����LN2���me�5˩Z	w��/�o}�?��B+���ð���~]�c¸��oh��8M77W���+�_���#/0��,{p;EI.�T��פ��Tٳ�`E� �&�2E_�0zPh�ޓYrh�G�~��%((�u����oO�tǢ�]K����ϩ��\�����EMMM�B�P�u��i��h�����B�F���uɡ�����m����Rj�p��ZǖnLf���������s��
�L(:���Xob?�p��p;�����v$�^��KMAA-�91�O(��G!���S�G��|0z���Zr"m�@2�~�5�#�R�__<���%hnE�K����D������x�$o-��((,,��tZ��p�T�+���/��Q}�+��t�oTq���}������j��x�@�H���Ov�w��`n��?B�fՍ��]ؔa�=A[�]/�|N96:��$l4���7�i��fbh�*-�'ϝ�(�W��;����{4vg��r���tJ�����;���š�̮����,6s��z�`U>Ö�g���4Vc�IS�f�㮖Q�F�B�@b�E��ZZ��Q!I��ǯ�dT�u4��G_#�0���;����7��p����r��K	S�. �fwV7kfǲBc�E:��1��O�Ạ�(�e���V�=������ʢ�e�(���k��mt߇ܸq#�襺�^����g�2g���`D�g}\\�f�L���~W�l�)�)���c����/x���P���>_�)��%��bhRnRt/��AD��vQ��Ɠ��琤��k?�m��4O����n�[U���T���Q�H\\�Lm��m��<$�i�/6G2�������;�u��S��^�����}��G�/k�m��=�
�^r��V��ID*`��H�0yv�2�Όc��bzF��7�\�9q�XnC���ɉQO#�O��
fc�^) �"�s;�B��3S3N3^�N�g�VF�����)Ge�-غ��dE�ۓF���h�[p ��Ǆ؋�p�,�{��p�qݺ��[)I���7D ����]M�����Ҧ�);XQ��k�@��� "�r�n���]Z�������V;��OE�[N�PCU�[����u���G#����M#�����c�E�t�F+�W9ͽCQ*�γ�atb!k%&�a��+t��"[!~�&�>��A-}��/��)>gI�;8����f'��Ѯ�}q���Q v��$���0��KDW��}t�b�wKWCS3�O�	��	F��f�au��*=��qG�};=���e�(�7�����P�����H#��߿�{���mG<K�(w���|�� ��zN�[���-ȉ�uܻ�[[ۆ-ez�����%���m>[���x���/*)�� G��Hw����[�AL5�lEaA�P"��>�U�T����B��6q�H��;p�����J���oW|ǒg=��ӗ�O'�"�{�	FtM�1��a����=��"(TC%�z��K���e��Pt�EsVCCc5��>Ĩ��B�h�.�&&�O�>UVV~J�J6��^�mTeO	sn�h|�D,i�W{�4?p!j�MP��,�wj�n��nl�5[��D����s7�>ߠ'��_:�fq�������I��+M(���Q|��_�O����i�*֯�xrY�W�8 ����������0� K�����*�$��Ǣ��Mj4�I�1����A�J�L@��J��g��k
�b?9;\o���>үq%,��>����]��ʵ�dd��rC��j+˵�H��)����[��c��s��t�<�[�؁��2r�|[��CUw�JvnnJ���E�r �1"��nu9��r�w��lj':�"DT�܁���V|���w��:d�2�{|�Zl���ߕt���B��_���5��!}���t�%�G֞�S٠W�饘��r��v��������]-���M��7�Kt=�tb��ʼk��0�Znt C�-Z&��q&+�����ћã�f2r��L�8OnXP$z�ih�6�u]�v���V����w]��kp��I3Z�~G�!�Y.Yتd��̡�P�e���9�����f�ܖ�[jw�j��)|�c@���t���[Ǎ`�T�b�z�k��?���q�bTS�^��J��qq�fЇ8$ ��{�?v�H�F����Vl SS7�C�x�$Zi���Bt��A��

�z�fe�*|耬�d8�%f��wg�
������ٞ�/C_�*������<A�2����{��pT �t���^lڞ���X1��11�l����k:�5�qr'+-��t��̰FrМi���[����w׵���`̳M��[��>AP�'k��s�$6��������M��9s��]G����7'���r+;���_���h@F��e�E��f<�=|�Σhh*'�����l���@��d�P3�Ѿ�k6hy�{��<�	�F�#�ڥtp`om 5�$%%����N?�=�Ӯ��-��4��yy����P6�ZZ��30_��/4����ǟ�j���l�.���k�e=���I>=aga�!V���d�˓*ș��ƈ��tq�����Z�x��a���1�>bfgW�=sWG-��ٲ��5K�.l��/X1��R賷l��T!'T�OCa��ʊ����C�zN�* 
�EcJ�W��S���/��#O��}F�E��.[@���=b #_|�9S��==��:�G�q�\�e�ۚ�\�/�!yw���L��H��_�%�#[ ���R��<��4�3�Xc����jbMlze������e�~�Z	rv�n�1��}odt$�x� �
A�$��p�:A�F������yW�3��3]��З����p���ĔX�q@L�L�L�˳��3�J�i�P��@���)��hj=7������{�+��4ħ��8�!����a���K��tw�o�[�w��������;�E�>�
��$0��Υ	<W]L'˭������E5I>�^_T?N�ݧ/!
������Y)1��?��~"����==�8M�P,�x�8m@�e^������х)o��Zb9)5(�6
��H��Z ��������,j�ӌ���PL���X�R
��d�i@~��(��Qvl�����g�5U~�ᧂ��@�H�UTz�i*�dg�\���lgI���^�<mm�/�vy�>�3.�9����ߡ}$��y�$3����+����[�}��'~Z�(p�ͧ�3{���K��j����� nzČ���[w�л
P�������ɂP�aw��v+!>Go��4���������L����D��5ow���+UU��Cau7��-d!����vN�Ñ;��Sp�p��>KuWW�ߋJ�8r��H���~}��Ӻ��˶@�8�Z��-�C@Pp��~�U���)�{�3���Ji"��7eԿ��҇'乭���)i� �}	i��ʘu[�g]0D&�x%���qqq	�:wnF���B_������⩨z�`�M�R�X�䚸ryg\'((p�k��^PP�p�ƿ���47+�'̠�8��2���̮��\��_��A��R�?め���4DYN��R^P'��{~:+��c�Cr��sՄ�ܛ��c�g`�u�پ䚟����á�"�� ����,|�>����˗�	S�W4�B�Z���/8|����ǫ�^a���o�+�r'�=����<L2`O(((�
D������/MLL䕔FA���el�-��t�JA�杏�?a�����B=P/ꨩ�Q �Q���Ų�xWśO@N,--��Mnzҿx��P��&p̊��#"�����X@�8��l*'�/n�MU^ڜ|��&"bp�Ν�����x-K������~�"��]������p;̜J�����X�5vI���F��������zz`T��JZ�����N�"��7�\v.�<s133˃G��y�-��ʺ�t���۷o��%�-^ך���R)Mn֛��ʽ��s#2�����/����/��{�"8�A���wt0�ǇfE� ��q�w@�`�/�O
+*��������a��X4�4�\�d��bXɹ�'fG�r�b�&��/�HROAm�tc�>\����c���co_d����5�fd�4���к�Y�d������fv�b�$$$9@N��RG���k��-{q����}�'�fbg?�󂓰����ï�,���RV�	`6���e^��13�*��P�?M -%L1������M7wVV���z[;;��6p�j�Y�AR�W����A������K?�7n����t)tv���!"#ˇ�1lДXC��U��g�������.$`LuD�uu-�OӰ��ϟC�}W�UUU3��-F����7��"��N'`�zxT@/zJ�����~UT��̈�|��u�^�.?��3�ŀ-�U2��Gg��<�w,ث����z1h�z9�y��F���e �.�E�*+k����V�C�{�����	2��߭x���_>�����>m��w� ��9�7Z?�u���F���k������Ù+�n��zg��m�?��������H7���B�]-��Z�"z�/4��wE��xk��DSI�|��$r�[49���u�.��Ȥ���fC�Z�i�*���0� O�^��<��z�n�Y���`xEPSo~'_�7L�4m��l�6w���lJRy�q\��%�e�A�R��~�o���/J�g�z��Du6e�%�PSco�n�ȕIQ����>�K�2>۲�e.���	gO��v�Ք���6
£�7�r���(�4}7m2�B�=#�!�ɸ�E�r!�?���ذ�-hvR���n���iZ��U�������Ԋjk���N��+/�B�tiI0���[<f��׿���WJ����FU�w�%cЭ�]�fl�g����n���9��z�Vx��7�%�geF��W-�`e���5�똯�!�3Kn��L�����E}��Q��Ǌ�4S��ū�������&E�k�ݿHv��G6o��i��a��u��
6���|����/�k���W�1�W�ή�!�p�h������q�\@לs����W�m*IS����hy'��8�K$~9L�>$���/x}�2��M��ɿc��@�dA���\M�a�!�*��gM^�x�������q�տ���Y�;�ߛ����L��t����㬤V�O4��#[�Ő���$��_o "u��$�#�-��3}-;w½��ѷ��w֜������yo�����uV^^�b���O\�weeՐ���"��.9>���$$4U�Xk����t�u�1�cʨ�����
3x���Vȑg��kkkjj���6'�8ڍ��`��D[h�'���������T׫�͞��֜v��?
KSը��[�t|D�cܩLE�u��]~q�&p��F��_�T+//wJefcs�b����KCO���ttTT|����E�E�&���(G��?����[�		�MM���,���k�x��0H �����xV*В���b�L��oT��#�y�������77t۬"���k�Ne�/�ʏ;�ux��޽�O7�#�*���SF1��}3ouu���^E���
L�x<�>�``����д��S`5]�ܪD��q+�=	�99Cf��!)��}ܪ"Н��,���U��-#ҝNWāXG:7~���D�G�"&&f2�!��c����S��%��!J0�}��ɁBy����ڭ�[XX��G�LO�~*�q.|��V�M�� hubOP�g�����bI��םT^?6.{*
���F��S�򟊣"�^{HEUL�����MB-{��8��gx�R��tL����߿�~H��z��P�S�b��t�2_�߁�t}7��d
d�ӛSu�b��GX`���@�lr�kv%Z	�敓�!| hNw�S���q%kh��dJ�տ�ל�v`|�Fk��$�z(>���u��Y�1��n(B�w����\��q��5؄���^~�xo�m0F�"A�J�`�e�]Op��a�z����{��F���(�}�s;VCU����ys� IVkN�}���ͳ|ֲ�}�a,������t띅�g�,:-�����k#r�	#)� 8vY�?_䈪q2�Z���%t:g�c``Xo	g	"5̋cѶ�V���6^�� &��R�f7�K|�]�;���~J�zϭ��Gi#�>)�����U�j�S�D��%XaO�)X�� ��I�u��	�L�<���Y��{�]����B4�!��M_��(���ʖ�����zZ�k��OV�cTDĈ�Y�V�rjԱ��^�#|��cc�5Bɷ���Ql���1)�Qa�0%��R�cn�i�3�n�(V�u��v<���U�|%HC�nڔ�3�nx��CH���f|` �@@�H�-vDf��[�������S���/ܞq��^Z�0>�}�䭮n���y��ﯬ��T�y*ד�Fx��������NZ���^GC�����ҏ������̜�u`7WK��Ʈ�=��{oJ�~)�����!~����]HH/��έF�0e�%s�i�M�gڱ�����ʂR�^����ݜ[�6�}3X(�E.�E���)q�yy~��¦�X���-�ݕW�Y"N���y-����˳��ͣ��U~�*E %�[zMS�='M�M�[��1"[(����RaZ֙/E��ZIKG��E����"?h[�\7P+��3�,=����N�x,�s������tx����ȱ5��]�%B6�/j�.��.��2��
�V���;�������X�)L����R��'��3��58��j�)NB~p̘��/�B�"����߮X
���m�hܫ�G��R��^� �r�H���ڏ0z�Np���r_�'+�#������u�GM��JF߿��}�Ņ�7���#4��ϲ\xHs����/?k{4�K�^���4��,:�T�]�/�����?�������o��6��f�����SW�@:��'��s�����S$�0]��{��M��H�R�P��ՂX�4�PU�&z^�� -��7�a_Cr��{�"pPzg�n)ߖ��kd1u���@�7����d��y�rX=i_w��7n[)�^����y(������J�XV���K�Q���:�e��$!�d��Ծ��o�%�j�2��5�K$k�,#&<66��R���yh���褣n��K`k[�8PSW�M��zQY�T����,��Ʀ#Y����0����re_nj�F�o�$�{c��
��#Go�
*j��}���/�쥴����ŗ�Ń��cy��������{��� LJBAEZ��D��[��[�P���e%�ZVE@�^j�e%��v�=���=������9�3�\�̜sW�=�k�մ[�)^����4�X=d����-�\���������"��^V�]��V���H��17p�90T=��IK)��"��*ƽKW�N�sRNs�.���r���딞<	�����A|�{����� ^�)F�b}�]6�j'�/�ʟۜ����\c��o��t��7;���.�cm�8\�SJ+��>B��Z��0�>��t
�At|�X;F�'T��?�*���Vݑ!mFݑ�"�,�>��y���*H��7eAp|��+�J�����*f����v$�}\�@iu�X�lU����jC��������`�"�I�D�;޿�tyR�<Z� ϗ��Run����������.�Xo���E���t�;\h=T\��b|%�qyɧ�����}X�o=��X��W�}3.�*�
 ��V��w��0c������]�e�{�9���}�<�I��.\X?�S-w�>�B���n�ƪF�b�7%��/*a�f���M;�U�6�A*q�"b���>]`~�tc���I�0Y�	����Ө&�󴝄�Z�R����v.������on���哪$����c�ܲ���9!.G�B�{�h:xQ���w-��jO��5n� �xT컘��e�=&�2��JإW�z5��h�%O�Ǐ�����ܑ����%�L~Z�0�tp��+R+ ��E�wJ4W�����/�W����f��wE�j�kV�PO��-x�����C�v����@գ��Æ�[���/
��w�v`ݓ��5p���_^j��<N�����=w��_����"�������U(�X��^|��1X+yS�u%��Q�>�0����ݻw{��Hd�bu��_�ÊWѸS*��b�ݧ���jۅM/����L�*a}fW��6Us *櫄Q���YO�n���|�B�XX��2]'*�ܱZ�Lr�:�Į����.P�vM��B1my�~H�l�~����irn`�S�UDF�^�x4]�������f�fЮ�ha�:w�\�������F	�ۅ8Xqq�����W4n��1~����O YF;���[�L-���*F<p�0o�%��&7�ۻ ���Z��5��2��A �ൌ������	����������hDv�)�7�$�m�-���4ظc�bk`c�ڄLc�� Y�_C+ۺݿւs:����i�r�|�<U]2;7{���v�-#�j�*��jXgg��4Qa��:�&ő^X�c�,RL���q~g�Έ�,�S���u�8E �uuc��}f�ћ�P�fɳ��^�RR�d	�����u�cNM�&���k#�������(���d����v�T����n�묩6g1[`C���p-�;��{���U�h�§�[+H�){؀m]Vsh����c�O{�VY-{WbF]/�h�Э)W�$HW�6�S�`�7@�R�[��aecc#�ةf|�]A#��}r�����9�� ��h\S�by�Se�E�G7y:a%EZf�#�
�I1Skckejډ�'뛈��L�1����n��ڎ,��i� �'x�Y�'"G��~P�>�ဈ��Y�z��O�����2���+�$�uY<�3��#Ѝb[����/%�c_��M^�|wS�>��q��2õ�"����C�@b=��8���/=�O�|���|h"Z<pc�7���I�<��{>J��=R���sG��� ��d�
�DI�^�O�ub��8��g7�j�=����׋Y�I �/\��jny���o��{��E���i�a��VvV��e�?�rh�_Jf{W��(Ֆo:�����sܼ�x)-�)D�X�e���Zր�����ى���p�"��"��.s���U����G {�%:���������T�׷�]_H0ʯs],�����}�:���R���.���x�����s=���wn{�|����=�����(,��Z/P1�C��(�C]�B%}��ԉ���'
C41`��%��x
߭ly�*|>Iq���D���WN��2OY�gN�tϒܕ�/_r5aA>�##Ï%Y" y\u�p~,i1���F�����렊��\�&^&�bH�k�B�+�߯���xAw�c��k-��Ө���ps{�ٹ9����(�@��7�Nfdm�&�;چ�D���>��~�(�R���5�V�l�~���w�wl�4g�V�����\i���Y
��	<G�|0k]q���gfp�ɖc�]�ç��W�Q��w�|Z�<�o:z>��}�������>��oX�.iz>i���T�������B����>��􌜩�t�G�R��xU����@��2�g֚������Z�q�.Pse��;��	��g���l�\���Sa�Z�:�Q)aލ9i>��� ����(�����1�,����ѩ7+R^plZ��|#�j�<''��ch�|+�U;�sy�m>4dw����q���ȟZ��'�qW��6�j��P���]C����$&��==Z:I����dF�Ic�GT#�B�*u�.�.Ph��&GK���tw�U�8�!m�Qđ,�ͷ���@Lދ��H�Ў���5�V��a���-�~ncccN�N�K�p��u�;�55�N��A˵%L٢��B;��smXt3��+ζT}�,!�R]w#`<}��o�s@�l�],�w�'LjZ�iKF:~~��:���v�Ip��O:J=fτ[?��J�����ҹ�㿪�-�ʺ̴2H���ub��$������'��rNR��N��l\�X�L�����o��B,�Z$o�~*FU}����h�@�F�65�æ3C�(J��=4 I����+M ��yn�%?|��h�QIi�``����Ǐ�Do�:h�ok{�Û��7�������;���>̖Zj�QsYG�t@5�{D�X��}U�@b5�=t�߳ M{&��x\�-�A�H��&�(;�94��Ĭ���dUUU���������?�8Fd���R�[�6�EvA�}H��H]:MY���y���eX�/L9�&�$_ܡ��[�:�dA�l)��VV��P1j7�p�8��UTV�0g߲�m�ĸl�2>tʬg�z
�tqa!԰��Y����{BA�t��#��T�$H
���Р;2�*ك1|Ĺ���#��%Ƣ��%)(��CL���Q�ШS�R�4�}��T�g�i`��Y��ǭyr����9h��;1kW۬�?(l�+�d��*J+:�]XX�F��������@��d���R
�'h�;��z/� �h��n��N��1����]&��ZWqp��.�N�Dฑ�`���χX���Y��GAaA�m���W�]�r�& 3b�ԟ56�pZ׹����6U��г���K�#wv�$R�~c�����gg�X�7�w��X$�4rʤ���x`��*�,����Ezj��xɆi
�����7��Ao��/mak&&&;���pIHL��E1=2�R��'�z�/#>>��Gt��M�ju5�cb�@Q79$Z�GLL�7a��a�#\�LF��N���������Iϩ��L7�hڗ��y"Q����rC?.i]p^N_c3��!O�Q��R�'N��uzm3`��9e�⁺�ĵ�q������K�}�H_���j�N�LC#.��W�٭G>Wv?��]��81k�(l�w/��ȹ���=���x�zo�z�E���X�Ҹ��l�+�#��䙙s�����?+Mklxt���:��y\v���Ѷ��2�ƛ�%/���*xԸ��%���*�ق��C+�����@w�����Ý�P*}a~���V!r1�J.N)K����6�v,�dhd$���"��W��Z5�u%a�g"�eZ���ˇ�\�$��������/Q�y�fܖ�׌ �.���ўg˿��� �[T �Y���ٳ{�8y������'j�H�Jˮ�_%r\RR�*�%e�ϡ��ql��
SY9��T������D�4���F+Ջlⅲm�bY�gC;�F��V�W/]�ߨW{w�f���m�o�&0�65rqś^1�g���O�N������#�&C� �b΢�� ��[�S���p��u��^�{46U�	���z�~���Z��p�҃��4��V���j;;��{����BB��03?����Ǘ#�7����K�mk��(K�?!���sM�!�N�0�����e-��Ζ)ф�3X�y/���$�4G�'�,{X����V�||J4�[_�=qZ�	y�{�� >A������׵��ߧ��tH�lj��S�-�6�V��U�F�&���'�"�z�5�S��&�]���'��	2��p��:G��u���b�;����n�����M푆��"�]�h��u��GVh�����Ǐnã�{Ҿ�뙰�I���NmT�xGG>C��v3���q�9p���2���V����1$e0�:���"%�՘i���hӧH΍�����N��{�:����<R�&����@}�a�4��[/gAj�ޞ�������q�V8�V�*�5�����ʄ	�0����h�ѭ��6��q��(�o��7�I�DݑW��]�,�B��N�]�����*v�ƭ��-�o�\����sj�@�3[�a�T���3�e���[ZZh�\{W
2���$��E�:�6�&��\\]#/P8�ꢐJ4��0r�fΏ��u��=�Æ.>�v�������e��q�$�KTt��/'�>�>y򤰙B�1�#��l����������Ӫ�h? ��S.��	s�W��I���^����*��4�������WH���[����yF���C����nP|�ߚ�Y^`t����f�I���,��T(�v��lW<c%���:�����@�g����qB��z��cm�9�
��(��{�0~N�vR�w>���zm�� �q�-D4����ڃ�b�t �Sܺ]�SyeRU��'�rU�l;�_R���6_+{��q� f�a��o�0�^_�2���%x]��X*v��@�J�d�{<q}�(���hg����oMO*qnp}�,�,��%e;�^�'c>�x�K/��Ȅ,uW�V����p<��SZ�mZ3�����E�uo�����c����ߝ�6
��e��u��E��3�c�W��e�O��z��Yz���[�N4�l�G1��J�V19�B�O���a{�SF��]�i&}����쇜����c�׶����w׷�p"���9+Z������ ���WgrB�'��c�Ͳb�ˡ�@{?���ĩ�֘����c��)�4Z�0��s��5�L�x��wo+��mt!�����8����sW���T���^���H/�8�23�[��hWC 9 jƷ��2X.�!�H�,� ;�E�6d�� A=��؊�Q����b7e$�Ř��F�H&S�-��
²c�H�c+}]��j*YC$䝘*��fo� jA�yu����e��Mw��i�K�;��t]�t�]�<t/r]�rW^�s����0V�.�h�˻>�`��A��EFI�|A��4����'Zl֛a�.�d�T��J�Id��I�:-����u_]{����Q���J6���1,am��;@���]�mP�4^��0��g���b���k����k�+�>�AK�|��5�^vf�����������_䞩2
{��n��p���M���5r�w�8i�aR�kH�6�+-{9�w��l���~�f[v6�#ïb� ��r��7�Vm#�E�쓈�%��5c��Q-���-z��~'~�������J��P�>!ꪡ�~��ϗ`�P�؝v}��Lq��xS�/n5CՄ�(-tY�gT\��ަ�"o��g��\���~h�2e�����
g�h�Nw/e���C>���6���by�d@z�e�P`G���N�n�V���Y.Ȕ�IS�>L�>�*;��>,@����wBǼ ��q��+b+�ؘ(�ʸ@&B�`�ϟ?W74,��re������������^U� 3u��$�䫂������������
�W�Z��������@��Bzz��Mu>(A=3N��8�!3#���O+7�V�q����~����ԩ��q!�U���ٍ;�bi�d�_3��u��G��`��ůs��C\�s\5*�� �|�$�0(�xP�iyz��I���/�N{I���y�,����#����ֽ���x�P<TZy�;��u���߻��Rs��SAPW+�s7U+Fϼ�P+.�q	�K_�����ɫ�rk3���������=��<3��\k�@�[ݣ�����3�?����"�5TU�������Sg*���h�\rkkB�;v<r���dW�~�%����-�b?�ز�EM��P(^HX��O���6��WZZ	�΂�! ��ӑI&�D�6%�/_r���:f����>ZR�j�!:V��;�$ǝ�|��,Sy�X�@՜�ӧ�ߡ�&�Qe�b؅��24�;�̑�A��$Ҕ�YS�� ���b斖���@�w~�Um= 'z�~�LsX�����)bab��g�G&���W��V�o���8�6�O0����~�д?�W<��);�}x�@����B*�8���|�44�_��Y�yu(��hYӢM�;4�%�Ѩ�����%���rr���M]�$6.��ZF�ݒ�����M4���b�����
�qP����M6�?�<֬PR�PzU�ĭ����+�=ǫ�$m=��MO,��Ľ�I�5^��IW��=�G�>}� U�T���CW�Ej�⤤w���we�!BG��)��0��f[r���2W�+����������a�%e\�,�Z?1|��
�3,��G�/�y���B�(b����8�#��I3PBx��]Z�8�Á k�	{b(�D�/e��*��E3g0ee��a,�	�:����qȂ����bPKj̇��4�Nu��r�K���p������m�f4pi��ߒ�_-d���O�ϼt�*ԹtN�0����A�N��7��y�l���y��a�3��b����Yɢ^*\�L��]]Jgk6+����ǩ�C�{��;ѭRD��X��{fC���.����n4����EF]L�
4b�����~1��A�G�����&/�]�Z2%� �~�\~jP�$^��ߢTlD���:=Li/B\��Wc}e����|�H������:�<���(�F�ՅE8���^r������t|.�T�Tem�ׯ����!�|gg�ۉ�o��+d���T9`u����1]�o n�Ǳ�ո�t����\���?[Z���Pu����Tn^��J5ow>� ���k����{�QD��'�,�I���C��2̯���`�b�(FI���p�L�K/���SN�;S|��Pm�4�)^q��/HD��߂&�~{V��'�B���NS�	'.����@gۚ��=6����/_Vݫ����f��!�b������Is��gmf�(��C*�YR`�����rQc��i��&���Ҋ�z�Zy�2a��B=�Cu�c�z7 ƛ{�{��Q_��N)W�fQ��X�SWW�4����+����Ա5��la�K��NeXu����3�x�t�@�y�Z!|����F�?�����)!q�>#l4*]�e�=�,�Ze������P~iR��*'�f��x��)����\��ЩW�.�Pv������ֈf��F��f�Ռϙ��!��n&4Ϩ����h}-gggw��艥�,�6Vu;�T^�������{9��r>Չ�C��s,Wt��,����G��n���'����Аm����'�e��c� �@v�����j�|!Nr%7�*++|v�e	��F�+UB��o�Tۃ��ea���U���K�N�zzk����)�g[pqs9�>�`���������xb��'j���>	 �z���"w$�oc�J�,X� m;�!��5_i�щћ3� *;'��W�i�ʵ�X&1>�̓���r� slq����� g;�`!T3t��gg9��[��)mC�g�L:�D>0��T`�.�Ǒe�����3�,ϒӤ �=}B�~���KMY݆ns�-M�F�[ ee�O�hjZꛅ��ʛ49�ϭ�R�VxWB���wJ�^��ZZ����=�:����뇚�b-��2����g�;Y�=���j7�'7*�ggg�`K�+����ᇴ�	��q���u��_,�D���<ë��$?���*'O�_�v��(���+�u��]s��W���9)��/��3�����+3�a�k'�����<����oJ�
y�4��W|�U'5%X�s�+_1en$�qPd��d3Tl�{��A�PW7�0��������cWr������;Al�;=�֭&Q�8�¼��w�G>C�A������Y�,��U�em^9���D_���l��_:���T���טcѕ\�{G��� ���}M�נ�Y]���J��.!nQ��v�i�_�$Хޮ���mR�R��~	Ȁbk��A���0%]βGX�4�#�j�����iq������'%��^g����/p9�
�zL��hi�j���\C�:�sm�K[�;o���罜*�+qJ��R�5a
>��/y����W~�ut�m�g_�zu�� 0�W�"/_6�k�(m-t@I��b��6����QoC�+޲o�.fj3뎹���FE4ڢ��9���5���-ù��e^��*��5a�*�����'�m���	�vF^���Q�$w�^ڰ|��?��#�%}�������p���[��{C�kCA�e�Pc�hMĔs؝ ��7[�e�VM��z�5A����9��O�۠w�S�i��OUU��G���u�:d�Si����Y�9r��W�^M�E0H.u����$e�@r(�+(3�_�8Z
���ǯ,�
:+-�>[;���G}�5G$)氾j��d��a��*��p =+s��uu����S1<xG�ꎤ��6dd�qM����g���Wi��8�<����5mX?t����c}�H���B|�߂z������TvSY��4���èb^NN��L'~kkk�%,?8 �~������6o�S�N�|�%���9�L~�b*W���?���bs�P\%��W}5}��b��A��b�Pc��/���ϵ`5�`Ǫ5����GkjK������0����[�
S�I��,�pHLB��N̗��2�}���w��"�MS�f�b��Eĩ)n�215mޚ:�%%�[��X-�М�Ä�Z�W���uJ�ǹ�y@�/��'�jo\�š�M ��Q$�j���e�����7N>+{�؟��u�顎�}�	\�GYi�,�D���z?U�ÝI����o�O�!�;3gX�o���W�X�;qzOb	Ҩ�4ҥh��xtGiϦ��m��C x/��{�,�J��?v�!]x�\�y����)QU+贩N���e���`�����,�荋wΦa��"�1��ܺ~W*Eڱ��������?Ohy����m�xo/�,�Z�;M%�1����V�P�m�c[����4[��d���vݮd�)��)N͘*�߯��O���Q�smk�K"���z��H���$��ƺQ�lW�Q�J���))>7�����42�s�(������ޠ�AG7bmnTI���{BC) �)_1���]2���%:K6,(��Q�hݵڮ�9����'P�j�����k�5]�Y�l��� �Ve���p���$�f��������~�I��!���!�k_�!g���ye��k�_���t������<q�66\ƒ�-�%��Q$v\6Q�9��~ۖd��fˍ��������빯�1K�i�y�&��h��׻�0
��&�����.�ހѭ�%Ts��W����U�����~�m.���Xf�[x\ ����pwhge`(K�L�܍�w��ۧ����klb�����
/}�`��q��U�)�����O5���.Jb����Ue*��(Ƭ9d;�����8��	�В7�v�u��>��n�����T֥�w�)��mNu+��&�e�X�[Rܯ�����+4��T��:��szx�ڵ����O#�@*�,����a�v�N ׻��x�Θ^�^�[$V3����dtj#���=\*��Xڴpz����ӑGj/�CTG����ٻ34å:������Y$
��je@� "�+��nҕs�ʸ��:��I���|�s/�PM;���H��z*��l��y�]������c�֭����͖ұ��k,!p���E����.Wk�ז
b�஬��<*��f�h+�A��ѵuC�a�b��BV��
�UUUWG;A	�ۋ��/iß�����s)�p��Ez�ȸ�]��@3'C)+�Fη�ՂSL|���5�����i�cu�N�ᾣ�����R��t�X��ZQ��o����+ �[P|�D�H]x�����Ze;�~�B����)W.vչZf���[�P�f~�j�Ѫ�Ck0�� ��YX2;;��軳�
3�.(������G�o���˘>4�C6��e�m��� t�۱�>�����=7�� ���ID(�x���sa�&�z
��F97%�"bbb�������zWu�a�Q-���ﶌ�2qrV�i��k�����vp!�W_fW�/ħ��_%{�L-,.ڸ��^��7"��C�kڎ
�B��u�~����x����9HDk��+s����t�E����8ڿgD,�(}utt��������Փg-��&tJ1�����{��N����/��6:V��6F�Z�53���i�JmE��/_���	@E}�
�.g^�K���V0R:���]W��1tk{+.)��Ǐ�7�j�6�G���;�:���F�Kz�I+� �B�]"U�,<|�d�HhecG8`wq��6���RX,�G(�pޣ�n"�C��%Z�O��R���r�I茼t��U�Tϡ�i8��	�����B6s]-k5&]�#�SB��]�r�m1��������y��~ɦ��;r���m�w
��VTV|i4~7z��T�M���/��8�a<�Y袂CӾE�X���>�J˰��H�.uUV32T�{6ArR�y� 7��m=��N+	�r�i���E2w�Zp��|�J㍉:l5lǙ�7G#�7�.��s����R*�o@x�a@�+$3��oq�`�A����n��W&	�J ��t
�ܽs�Γ������s��uFK��Z���g!�e?�Xצ�2�[��{J�q�_��g��ԅ��T���ܐ�h��hip�XWDd��W���}6ȅ���1�8䖏�胋P�@��gZi���4�%ߣQZESw�k�����,X�!S|�#5z�ޛ"�=R����r�F�|���-,��N��ӡ~�N����H��??���US�����k�����h|�[�x������B��g\[U�}��������1��چi�l4-9`<��R�F�¿�)�!���F���}.�rv&*��⟰��;N��������쾊�#��+�>�S�d^�ɏ�MI?�p����0����N��Z*ҭ}v���Ҙ�Ib��� ">^i��V�?��@3O0�R=��6��Y�L�ɣ��� �{tW�|���1z��p���G�97���T��
F�}ݫ��v����mr
�;��_�/A�IXFTT4��_F� /z��)���|=����񧾀���T
��1�\��X��(�\���<��K��Co��Oui�>[
̒.�2���=���K0���N�|-s2��_i��]Հk���p�?4SA�A��j��x�����z�wb ����D��6��|+����=?�����J�\�F�=��%qE�~��Nk��|<"�Pw�g�<	Cj�?FF�Zo�H�X�J�|w���$Y�������<�\4�~�ڀ�ٛ	3�$R�Ac��E�#������x-=�p�2uK�vP��D����&�B�&I��tTn�-�u��`���2���a�

�E�Ƙ��`�*k`�N���ʑ����=29p�<a_���� ��w��t,mۢ�`�9�%�	��3�l_RS�<>=/��|%��8z�"�$��ߋ5���,G�����g�S�D�L�_#`#��v�w9�G�]����P�u�e�T��*�/{��jr��Y��'+�n�"z�����
7�4�5��Qx��8���|�"��V}�*���`��#M��{42�M�!j0D.��g�����?N���ԃ�~�G��GP�r�����>1����D{4�'�{n�O�^��w�R�>���r��AG��l���^m�5�O�%�[p��z�Wﰘ�=x�b}<CoCH�AT׺��i�����w��9��a���k�{.��m~�tW�e�uvL���?��We����_�L�u|o>�`h�mm�[<���v�%I㆓#��!2**�'�2���{��e֡H��e�.>\]��V^y��=hK7�w�`�6�}��5%���L�̨gr,�ZY�1��=kq����)�5B��E<J'�y���ږ�E&�b=즲 ���P|�@Oy5+`�/L�C�.�>�3t�^po�T���*d�`׶�TCC3��M���!mF?& �I����Pb�, �k�N�p��-����7��	����o`����� b��&1��:Ԇ����h���qO����_aJRf�_��G/�PRJ_��b�ԭuz*J-w�S���e�ip�ƚW/ugA{'��K��'�<�?�3S��/�j��Z�|�1Q�4��V*��� ����A/'�
i��j���vm��FIl=!��r�7rE+,���(�����A@�M柍b�����T��NcK������y����� `A*ʨƭ��ߋ,��s�@�ُ��Q\��zX�K?I���{6�f�t���{����SL��>�M^�}�T}>�{�((�57�
����uXh��m�w_"f��^����B��6QÎ��������J��U��>�H�O���b�_Z,z�7	�%��啕�U���\����a*4�HN�E777}�~s�U��SQD��_/#T�*(]QYY������օ��qh��Qe���Yw��.|��7�#/e�։�M�C�{F������ �p�d���E�[������:�_���PL����
J�][�?��"�n�¥/�4���m��rw0P{��3{u�~�G<(a3_<�}A��U��HN9�hE$�<QL�R��$%� b�`ѕ�g�"a_� ض~aXO�%���$~ݳ�ّ���D����س��8��`�qo]TLٙ��|��܋M��ń��D���X@>2WVV���z
R��mo��j�����f�ٴٓ�x�[V��V,���>Y����dZѮɪ���YGw�ir;*{�`X�>ǜX��׌��g�+��rq=G��=�nX��,��9�t-f��|Ui�uĥ�0�z"z�)�t�o�L�L^��F[�/�A�R��F��{o�h�[��cx�k�Y�%���**K����ju�mG����G�}�CZ��ۋo��a>a2C�L��63��;/��`儮b+PJ댜��
x��D����z�%V��j�ݡ2bhh�V�.BS>A�Q1x^�qxF1T�g�zA�A�Az�#m���6O���rE��`�]�<tI��K��=V�֑�4�;A��@����GVC���Z��y=sZ<FYȢ��/��fD��C`4w_�޾}[c���j=ԾrQ���|��l��6�(t�)1���w �w�HZ�e�P��)�8�H� �9�}JA�������K�j ��Ǯ�Z,�H�����X�&g������8����l�&�-O�`��P$�<#���Y��QQ��'������n񀮺���������x���������5����zDX%P�	�3�׺Ώ���\q�����,jj�h��:������kNR	�ͷ�4q�34,��rq�@��\���'�(2�$6��ம΍*]���Qo��U�Nh/��8�J�>u�,v���e1�d��s��r����>����^���w�"X��A�*I*�l�r�Q��C+����c��r��g�^����k�PL3(�~��6�4&��͍bw��o�
���*��D<�B�Ϳ�h�ݤ3?�������ܱ�Ŭ�Жz�5��1���S�����L���R�z7o��V¯pdX�b���e�&��Z*�\��ٷݬ!���n�ݟtt�1�4kY�ь<򠝛��]J+R^�A1�Q�����_�H��Y���R7HUqB�$?�Փ�O�g�Sg�F�J����3�����)�L�bY�΋fi��F�|A�������6�ϸ]�V��ʤԈb�j_*��8f�N�/⺸&_BG�&� �3e�Ŕ©kD?P��I�x���<%�eꚚ�u��.Ȟ��|��!f]J�����#��3����5�u�����/����Ӆ�ۧ�o��3qÎ+�G�b�T����𜋫���a�d��m���'�4.I^�#� +^��j����[��L�!ʠz���pF+y���^�����W��-����a���>��?(�18%�Og裪�"�� JUhC�V{��n[����&���v�\��cn��#��UΝ����cyg��t��[0?�j�-7mk7�X��0?_�_5���*��d������T���_k4T����6�6D���2�GM�*Gx��ǧX���W}}?mI~�Ь�	����BEqxT����'�Pӵ<����T��ٹ�kz�d�%(ر���e*~x54�B��X�kBϜ,/ƥ����Y��C/�Nwe���Om��_�)=h����n����������@��H�,վ4h�Y���M_Ǳ-R��5<??��>���S3���,�1�C��ܼ��5����}%�2� ���~K`�eO��������C��'����7d�p�M�M�㧩^-�]����H}8x����~��_�xttt@)��OIL̬'�l{a�� ;���Y���ocT������H�-��9����ffh��k��`PM�T�c�8��C�K{�"��Ze����t��*��ޛ����bb��a�0hz�Ҳ��3��T���s�5�n���5�B���R��Q��GǖLXcd�؍f	) �_()oεA�2'��L_�?ۿ=PhP��w�1R+E��������o��i4z9����q� /L�)�h�<Ͻ�L�0XX8��XZ�:X�#2�'j%�3���{&3���liY�
HX�i+QJ�h뛨�>������
��q����Y����%=�&��d�����E�g4��M���:�sO9�p� �������H��.�57C�b������ u�8-gɳ�wY��"k�TIKJ�*�,/>�Y��_2T,��^>d�y���P����=�n�����$"ު��T�t4+m���aA�G��)ɑuz�&��s[DiR�ss�9�j�����Ȯ�OH}�ׄ�Bmp�j9�����SY������B��7��w*٧Q�O~a� W��j��f {!�֫�|Opy���*�����F����l���f�^iz2�c��uެ�4�L7i!�^:W8V]B`�e��g�����xy�JM��իV+�y]� y������P���>T����~?^��B� 8�Y+�Zk ,�"��0��G`�G�a���7@P�{;�H��T�Uzj{��}ŖÃ�¦Wg�rF! n�:@8�;�+Ҹ^.��_�q�-a��Cvڨ��� ���n��l�q�+E���>�n�qD:���nr�M;�Z��B�?�tp���r����� uf)/�z^�ؿ���w��׻�3�YJ���-��=>q5;x~�%�����E\�D�����5�Seu�d�?~Qm؁����2�>~| .���8��h�</����~����n^'�	��B9���ǻ�(i��j�����ȧ�����:V�|ɥޏE/�.������Κ�^BO����Uh�d��r�/���: ���1ٓ%� ��tu׉�����S���j�ό�tz,���:�Fk4�|�*3��9��j��ϯB&�Ӓ��/%����u����.mDj�ДH�������y���/l!�]#��,�V��X��X��3g�7�H_[�շ�T:��`�a���t>�St�z}P�q�4��s��\7���a+Ia+�m�Z�rlz<m�ԅ8X!�~Sz)�T�����7�t�n�{��?��9>�NT{J��W߹��J�nb���.�؄���P��k�A��v�鐙	�6�4i��p���U�:{������Z%��6�6z�mx�9��qJ���j���g�C[s�E��H9��e�*'�$:Mo	�o���{�ѯv�2�k�ðk����^��+ዸ+�;��Y�Ǻ��+��Ȥ����8����5�@�J~ˈd�v�8���/�P�����(�\y��੷��cnii��O����{f2K�����,���bn�kĝ�.�Nh#~�[.�ke�����P�s�e�� �+�`��嫪�J�_�=�����O��}���:Ѻ|������Hf�#C�Wa�_H~B�cn@t��	�I�(�[0]s]��{;�M�%�F��)Y�d��k:j��*�5�F$���*P$X?�w.��.I��.�|#��ť3�j��Y#����р�ٍ����/��+�?t����|Ŵ����3�������|ԝ67�������
2-ny���`���u���W�/��r_����NBAA���hs�����;�1���=#�S��[��d)�|d"3���=�VnI^���K�����=w�g_�	趈�,��@�"��m���v�,W�g����PU�0�4r�x��J�c}�x����䚵�x��?�կP��\`bb�T��o�%)^�I������3���`��a��x�k�\$�N�CB�|�_G����U�YGL'N��ŋ�ѥt�U�j\/��ṭ�;+wEEG�~��(ƴ��2⍟e�Ũӆ���[���8?}1:���+ ����!<��NQo�g���Y�S|���+�,a�+��J.��{��j���5�ī`�����˗�M��E�6���^ĚaD����~cEe%t���
���v8�M˄�<�0Ub�Yl�J_��s`UV��h�-
��z��q,�ؘz�b�p��PcH[DLl�_YE��>kLB�����Ǒ�X�Z�]]q�M���JJ�E����N�3kG������^����#���ں��F�ѓ � z%щ^F	�轌2j		ѣ�:����DD���F�1|g�����w���$����Z�Yϳ��k{�>�i�����rp3\�CMM���(v\�V�$}Shi:,�Ǝq	h?R�,a����<@�w+��˞^~�Y��y�u�c}�8|3����"�������&��u��b�����EBڙ�[��&���6��q�0�
u M�������OK��d���)�E:S����������H��T���T�rn$���&3������A��r'_2�f�;����E@	ol��i��H*?�ϵ�8<c�C@�Q^"�r�e��� /mO��լr)��T�>��K��cb*��F� ��iF��b3˨��$ٿ7�l�>O��(����e�"��){�8��u
g̘;7&oʝ����Өes�FE�I�<$�[�?VQ�ˆ�ݕE#KF0��Ύ��ܥ��J��ٖU� � [�@5���1�~���9r��x����WZ��3�5Q�����3|�j�����>��,u������Z��q�B��d�\�ݬ�]3��-���x��kxs����!k�U�P���hy�����F�п-u���~�)옱IS�Qhm�6n�@y��n$�8� Y��v�&HO/ �'/��]���c���w`)g�ʉ��i���Κ=����2��mZ?��� �������i@Df�2���Ӏ;ry��z���$g�X���-�W��:"�h#�&?ߙ�������;K�}*�%���خ9��F�9`c��ژ[�� �Gt�<��,���jp�[�:B�bW	6�&��������"�Z�����U��r�	�[OB��	NǛ�%٦�l�������V����,O��	W��u�W�S���v�X=_�UsLYe���i�/}2���j3�+�UW��лL:f�Ժ=�dՠ�����z������b�!���:cG��5��೏P��~�a3 ���.Vb;@Ѱ��ү`������b��ť���:���ve�����]7N�3ڞpl�+K.�sZ������rle�cڱGH�ja�H5�z�f՝����Dӊd����>w �� �hkk�T��r6�`g��|*�w�&D����l���O��r��񟞤��PZ_�+X����!d+ۂ����Aɉ��r4BD"����u@{�'����D�k� ���.F�HA>2����#�wL���fL����2!6eRP����b/�gܸ���J`����W?����F�p�/C�=����o��-W�!6�ӗP�p-L��UW;9�w�LG��ГXXl�W�F���wܢ��'�li�6{���Ue�욫ty�yi����0'vu���*AVzF@"��L�|.�^|�_O)�b�.
��ֱ/�@*��ꪏ�;�/-�������D��`�3C{ŎP�:U7��������ғ��yv)�9T�/��~1��p��Q� �o@W�Q������L]�C�g�˥u��{�����:y�Z[��MA6��??;�-~O�	�o�xC��|Wu���fZ����h\0��r;Gެ����� eJ:?o�o[���r��5FFGo�@)��}F�{���9�����/��բi��N�	R>X�K�TD�t�� ����⺳M��O��Awc�_dOW��~�1x#����2B[��E�	�RM鞤b|/�^'�v�4��y!�n� E���	����t^F:�D��;`���)�=�'��6r1�ɘ�
5ߕ-��\7���%��}z�����]C��s.�2�@�:"�R��U��J��g5��������1R��s>���~;�����;uq��������C�X5h�1P�g�IE����X�>@P;#O�h�7sŉ�IT~6�)]�?y���Z�1�Il��n�����e�_H�=��k��Baς����u(��R�`�~r���֫�����j盓�c(.���B��>~���Eb(���8�(����!� ��O�j�Z� ����"� �_=���G��Fyl6�L�Uz�R�F6��M����͗+���j!2��
2��#��u�����S'~�_?-��q3�qӕ@���^�]�|<�G�&]
�C�WG�P��@��Bb����Pc�Zm:
"u�[�~����8o���t�$�b�![_H��-�!z�=�H����\��l�U�`"9���m/�4�E�!y���i�3i�;<
6��y�ɛKy`\����Zfz���@���mƢ��{N�/8��~�H�3��1!�b�����%dMz���+ש�*1͔2z8�@g�����B�~ҽ�Y��s�#N�_�f�Y�6xf���r?o�ȫT�K79�ټ�l(�c.`\�f	=msM�Oz0[MbD�.wa@mu�K%�ѫ{A5�L_�ѣ��ӗH_o=$�lZ�ʅ]�k+�s���N�_�#<���f'���P��|)Mg^��}/�@·C�a�<A��Uf��0��[E��~�Y�7��Q��L��po���wh}��3�:�-.H� �u���%���9�;�0W�u'NG��
��c���l}�|�6 >�'d)��?�L
�l>2sd����3���V��r�L��/i=j��z���+e����R|w���X�؉��K@'����u �/Ǹ�!Y�:�A�����'�a�l��}�#�ԙ�>�T1����3�e?���9��h�}ޟ�FW��J*�3�[��	�G������̣����ʹ$,��'�TD�x�Z�9Ƀ:d��zZkNj�d&��^����#��<�z� n�Of�'�]�]��M�D`AC��i�a�:جx�P�q�to6��y|)�B���f�Xض����q�q��G4��Ia>�P�����Hڅr��,V�K���$�vV�F+=A�m��oX	�Tn%����2a�b�K�hW�����E�� JȄ�o����!�O��=C=<=��GSJ�m<y:���##��:�dw:sOw�� G�Yq)X��Y�Y���>��5
t��mZ���Mm�y�`�JL���QJ{gδ=H/z��~��N�0��z�7K��d��:[(�*�Aq1�p�3]�D�g�|�1��?�ЬY�յ�u_��_7��H��Ɣ����
�d!��ۡK�L�{��iKA�M�غn�p{���7��Cْ�ly�;b�a�9�Ǖ�����յ�H�9�ѫ.�Υ�1���yw��@X�c��0�}k��Ņw�Kh�QK��N8��y�ǑM�0&'za�k:�e)u4�5Zo����*/"���ĉ󚫘]���h�~�F����-��;Z	�쿟��� �ˬn�˽;7;�yGH�o��JD���Rqܾ]�О  o��?Nf�����`��I��T������/���)��	ɵd`
�o'W�ˬZ�{D�N,�N��Q��r��H���Ɔz�ho��?fo!�/�=�V��ǽ��6��r���t��"�߯k��t5�f�s�p���$HX�m<��j�S�a<���.Ǣ`y`Xa�)(Y���C:�[��$�o���V�s\����{���/N�r�`���31xnP0�{�~V;�u�Sv���<�t�a��-�tMY^�鮋���e�K-���s�F�7�����x�Ʊ�jҗ�*�.���
Jj��F��0T
;�à����x�6�t�SEE�����1��ưHb����ς�t������]�2]���m�k8�[8�7��e�O�Yug��yʘi=;��bG�:d��U���+n?�'@"�e(�"�$/�q��ʧ�Δx�ୋ?-��j�g�S�<��lӊ �;�f�,qD�+���Н-oUg��*ፑ����]��ט����{�W�}�sfF�|�������$�s���!�
;83hV�*y����s��c��s|�S��sN�2���0#p�tk����W�#��tq�X_� �}���DT^�8��H/���{=��7�%���I�z{�XT��=�}�����E/6_}��k�Ԅ=N5����������&N�A�><�>��']Cj�V[LWb�
5S@n��TZ�\D�-�7�V�_�n�,[�Vb��_e���l{;<��񐃋Ke��O�-7���a���-L�qeJm�陭u"��붮.A�G?�Y�V���wY%�<�1�W?:$ZGo!������pΕ����:.�����IU���̖M�2������s�&tl�."xM0��	�*�3R'H�|�Ukd؍��mA>�(���Z����gT����F�|��3lK�O.h�
��k �\:���|j�SR�v��^���B�ԗ@��������]͡�-�4��5���ԯX��J�����4X�-ɂ~�#/���9x4Tb���
���v׸FP@"�g���6�,��G���)E��#��Md!���<;S�uY�ʨ�^���K4�5��٦�)���ڴ>�p���ʼ�F�?X��ƅ8��9P��ߣ�Ppwwϋt�C�ns4m�G�N�.�Ү�����Ė��������ܒ<ju>k�>BM���<����׋���y�{�C)hhh�.��tP�_�tiλ�h\]X��d�D�W8ߙ�<4^\R/�xp9�]B���͜�j�P��O�@-�+�Y�Kx��J�t�O��Hs���o����$1h��W�b�mo{UX���M@Vk�k=m+r>?���qO��;G{�z�LO[��봒.3��o{�.���Hr($UD7|����\(���龗G��"���b#h���wm�xv�?y�,�I���q�Pl9��~l��ִ�[�:BL��	}q�ی�R֠�/���]*�[E9W���wʹ_�8Rn]f�5rX����d�q�r��*��_�����NN%Iz��RSI�u�9��RA���21P�4�VbP4GoP)՞/�Y�]V��QF+�c2G5ʱ8�� ,R�f��*�@F�_��$�/�V�F8�n�m^7��W;�_���z/)5Z>Ɠ(����^ĸLYn�-(�Vu�o3�����jK'a��)X*��N�/�C�vm�89��Zi�ԍ~M^P�����=8d�6a�矬���:��rqю��	ЀJ�K��F@V�	
j��/�fC�5S ���	U���x��$����8��֕Í��r �}��Y�2�Z.��
��'�]z?G0#W��ۆj׭���ƊOH�7����n��6p��q^��^�ۄ���T��c�����VUE�r�z���
��N���n����G�c�W���]�1��� ��ˇ��}�ӎ\'�ãD�A�׉��a��dm_*��HŠ��3�-�8�e� ������xM�^��'n_c#~��QH�:c3�t3�M�[ZZ�%%��???e�uk�bZ�Q\��L$�D�f.e�Pe�3K��}�٭�㝈��������q��D��Z��:��^a���>��'v���|�R�o?�qG����ӭ����s���9�1��J�ُ+�ô�_���hy�sv�����x�ܓ��tL>]ʿض;����3�8���~���� -I��~���|O�z��!�\�gG�m7�����m�	�f��Q����h��qz�Yp��T��������>�9F|���4�E��B{�5�1��0�9Թ��!���s饱a�ǂ�*�W��7����'	B��f;�ʙ3gF��S�����⮑�c�Q�������ǥ���ǟ�8����pIK��.z�����נ�m0e	�J��� �~�F�O�?.s�>�T�)ڕQXyy�U�mv�]hhڜ.���D��M���-Xg��V��&]�Q�et�ː��!��u��K�(��f�ޞ1fL/_�u�����U����j}t�HQ�ESI789i ���X\�a&��,yc<-8��mn�<Qo����i?��~&��=Q�:�тi�ı#��X�C�K�b3^ߖ-�h����;M�cD����K�Pf$�C�l�����\�U�mŻ��'��}�U�;��T��|M���&�u�.>d4�dCF�?-m�d[�fY���"!��%�Vrq�`o�tC�zld �R|�m�g��>������=�_(�QE�_�u-�2ǚ��E/�p,X����U���&��"����6OF���{��،̈�1��]�����堽z��QE��Hf�t&���O*OM���'%=|�5�����Ȧ�c鐏V��$�d��� d�g����Lnh���N�5�8�Μ|ŝ�}�NM���Fh�ЋR��	�!�jê��:L1�N�E䎾�=�R���WN�(ww�����d|�����̭O�:|?�)��1����{A�X������-ۜK��[���HMc�~�d�:�4�UE��uwqj�o���<�Iʢ��_�c�Ν�[Ge^m�,i����}��Hs�Hs���J��H��2�ˁ�g���u��BI�UTԝCUC��l������A�`����1f���`*�*�[��@B�j�&r)��A�_�6Ǆ�"fjD�{���xrEJ��0O����x��~a?�{���B�^DI��j���ZG���GJB��r��>��y�I2g�{�K<3����.c�15e"�/dm�)i�EV�3�{y��;����m��4�W3dQ���:����d�`8�ٻ��6���!�����|�٫b5QE3���O�I�@�>�O����5>5[��Z�ؗ���XjET�f��Ï�2ߗ����98D�8B�/�L�v�/�.g�����5�<S	m� �)X��ɟ��x�fʹ�6�܅{l���l�/!F�t�)�3�lD3�4�q�Z�!1 Y����=�5PupH#���qحI��y}�y)��(� �C�Y��\u�t�D{�ã�~���(?��N'Wڷ���[�s��JU�F1]95�8�������27���G�U��,�(�B@wҶ�Y��?�Wh
@SPCqq���t�!3�oy���������϶2���c,r�[�bD�]�������56;l8�a��\ـ]ԳJ?V�N�W�ܕ���i��+�R0��� ׌i�h�t)�j9��#t~�D�kR~QFG��tHq����U�E�
YjI���������q$�QWo�������K�<��Svo����Z�>�aѧ(5��S�,�\��l:/-��iP�xR]�����to'�C���^K?��,�Hn�l�{���xǠ|�Xt:�e���-_I�:�2�$�gt6�������C�]�0�j�ēw��t����Zwr���m��cG~���[�j�d)�t�.����o��+~]r�1Ϊͭ6�jnL����#�k���Xkn���G9e��W6��<<ʻ,��uK���|�fG���g���&K��q	������p���"�$�&t����nRl,e.���bG^_��7K]͘�	�7��.�قNc��m餿�����L65�cI7w�I���3k�p O#<�<@o;��@dD�D�0��d����`R�F��r��.�~�W���h�x&�9{f�2��F�������O�ir�V�� ��=H>�Y;�}�"D�TGW7&T���/����t�8p�n�l�h���U7x'>4Y��%�_Љ�ED�ubQN["�Fv����k%��<M�oտ@1Ǆ_5=�s�f@"R���VY��kz!ɿ���!9%�C��,7F>��]��xA�+U�"ό�Y$��r��ּ|b�����^����@�#:±]�n��/��z�ω�Io�C�/E�
6�/����Ѫ��e�� V�c��j.�;��4�,WEe�}�-i��+�w�ܾm�b���{r���VĻS�o	��>�j=�»Tt>1<D��F���e��������;��OVUS�]�h���"1?l5 7o���/���kFɦ��_Z~x�|r���f�:+�Õ��8���t�x�	�j��15nq���K��e#+��jx4A;V�ߛ��&�G�/��O�hȒ;��x�����h�0��0��7>9�3�Nءi���IQ�$�җ37����>�H�y��Z��x0�c����B����\���sA���!	�-E�X��(�u��Q�j�0"��2�jR=p��&l�g%륿��bm�e��������
����	|��_`�P�Jd��cծC��W������|�a��_c)�v��S��i�\I[��Y֡,�s�?n&�s�Ҹq������vTk_a���k��?�aU�����e_F-�ņR0�O��.�}�h��y�q�ޚ�C:����9��f+��w�R���Gˎ}���Y�E�;��NkM����֠~� "or� �S�\�E]'P%����sZ߹��Jn�е������u+��4�5ռ�<��F����s�n�|��'��h@�D�Y.��W�.�A[Y���}�&�dh"��E���ݘq��k���c�V����*g$���yɪ��rT[�8*H���<��-�8�ɴ���3�s�Q�7M}�5���#�̖f�V�<��������D����dpWW��U7���}(�ၳ#��%~�Sj��̇����^�8A��G��+W5����;�Ga;L�F��S)C�zT�mb�%��K�.�?e}���E���NcDQ#��whђ��>�:�fu�P�l�;������H��m��d�ٕ�C�VF���.�d�e�)<xd��$~���Fi�ih�R�vx!>]�0p�p�>ki�i�X�_��rr�E�ބ���y>_:�]U7��A�q�4��o!��v���c��j�G���ud$�J��󸜊���(Rmc�N�w �(赂<^��"2Hg�4�X8��^�/���s^kK��/�A��m�?�zL����kYû(�ή�ޙ	���'`������M|wbP�"����R�����7� ���%�MB������(g�3^S*�g��>�����Z^=y��b! �����Г�*���/�8x8�Si㔬+�C
�?��~��]:� !�՛����p��9v�9��P�T�]���-*��L�}������J�#�!yQ�r>ٱt�;c|bb��h|�̾!Ԡ����z������&7��2]�J߇F�}E��ժe&[ԝ(>4�$Vr����xA]�[�#��z��w}�t,�|D����L5�0��z��X����[���7��y����k�	VRN���Z%���|'d%��mX���2��4�פ�3g(���]�h����555g$"s^�8	3�6;
�� �]xq	�%ZZ�}ߨ�D�0G����l�����#�{c9(��>@3����%&h&�����r4������wk�}�,����ic{��/����R-�X��k@/	���	�U��L��ďDwC�s��.o�i���;�6$�u�^�P9�:�\�>��\�ߎ����i9�]ψ��G�`d��B�W��O��Yڭ�yyKyF�C���x0��G���w@����d�{xHC[[j��Y���0 B���uץ-k�G����EkCw������\�� x� ����<�
~�l�bɌ�f��Ī�8�;��
	e��R&��C����׫x�S#D\2;E����L[9��پל{ת�h�In��]��n�v�J�0v�(�T��!��o���a�z�u�O�Y4q���,�W�l�h&�C��w��.���X�� ��RF~��P�	�1�ߡrq/��nWz�[-Y�b���u쇍M>qZb������Q�?�l�=��k�k�z��s��Es��d}��q�����*={k��NS�^0����v����k��aCٽ*����EƛR$��3���H�dv���6܂Qeʭf�H��35s�5���'��֤gX�+�K�(��|�&zC^˚�����W)��g�v��/�Mv^.�/��1:8"N&z��1Q��W��Q�R^H�Tia���y�*l$�5:d�����<L���O��p��b�܈��������wBϠ٪^�������Ya��'���-��}��B�k�>���� 2�u�T���`����l��X1�oN����m�����շi�$�^r
�܄;;��nGN6���$��ƻyqm�^�Y,�m19SA�����:֕9��5�3&��Y�+ �ﴎ�Õ?*�=|�{s�Ņ�Z��H��m@���<�x~��$�����T�r��Cf�k�G��.�m��X�NT.�2�!�����Ȼ��Z�|M��A-s`_����:��z���WM�ȅ��iz�rgR��ח�9�V����> |��œ�$�3�^�n�R�E+����g׿�L��P�[3e�g��j5utt���_X��cŇx�� J�O��ݒ)N��	k �I��Lr�_�#����2H#�� .�s�UŮ�3
R(}�����Ύ�~�����Ł���\y����2㢣�gv�Μ)..5��,.f���ődǅ�/:�.�	��+�Mb�j>�Ӈ�[�W��sk[Y�R�odߩ!��H�j΀�K4C��7�-
�!,��ޢ%��:	�?��<�_�$5}��;�2w�!4�����t����s@-GC|��R���斫fL���/}�����
���;���]����"���N��`t���ւ��Ί}�*Yf������BD��OR�����70��z���aÏ����~�-��|��#�w���0�ٞk�A�K�O�����z�*t�h]�-�圛��Gj��qss'�"{ӵ[J�2猌R�g�PAb7}g��Ƞ,�Mu9~���?^���У�|Y��#���R�ȩ��FMӱ�;.]+⪚k�}2��kM�k]�C͔2%�:�O�oIޣ���F�D�w!rB���z�8�[�!�8!+靏_�W��3ͥh��n�<��J�e�������� �_Dv
��ym��#��@��mq�$��";��ؠ��t�У��������E֦��O�Qۏ��&}��P�&�Aa9�+���с
�r���.�&�ޫ��tcNEj�Y���;�*�EMO�{:���l�;v���S�~�Q�%m�քowpJ�8�� �f�$:{O��N`�3���###�~����z`y�T�"�ƌb.$ޓ��T49�!	���ڵ�� 9�	Y��Cs�Ԏ��SC�7Դ>U<��IO�e�x���+R�� �>r����,	&n�[cכ\J`J�3 75��Pq���|Mgj�V�W�M�� ���f�z�^��#s��O&5�b	X���@��Cps�i����5�/�i����,���,iP�x�2�	T��4摅�T����NrH��L&��tU���_���hL��}@A��������ؒ�nҍ`)��w�F�(6s�����U�A��y�\K9?F�.d�[XI@�4�i�"]�t���G�ǍT�Yu$Iqv韔�JZ
�K��@�f���_�����{9[��$W��c�m�gt�ҿ����~���RX�QB^Az�N���P�mr��F�K�tW ��g6�)�]�;Z�����!�1�*���R'T�4�7��2A���Yf����U4�x��-EH��ڲ29�rnboa�ǅ�qii���;��H7ɣ�;M�t�q�+͸ޮl�#�v�i9����=*��AX�[:�}��a=��wX��x���rK��x�U��v��H#���L��!�Хn)x�?^ԟB�A��t�Z3x�*�����<<4�Ę��ٛ����lP!Yo�,#�7�1C�!����?���O�0
���f�6�j������
 sO0�C�p|||^I���R�b�^�W=퓑3]�"���u^v/�N6T��S0<P���e�=b~���eoAf�F��ۢ�,/�bV�V5�T�p��%J��xV���b���������ޮQ�؉���d)�k�Z�+#��O℺zw^!N�%aR��K��,�]=n�\�,�gB�]Nza۾�vє�x�2jk/ 9���}�k&��!�22�_�q>����Yc\�ɔ�(����7V��E�N"���Ve���{���\r;E�:��ijb�	����7X��5�N#��8t��&%be�ߘ����i������"�{kb��C�gY}~|��KNf�t�-���r~G�f<Osz��w/G&-�z6@�^�'��UD|	�c���I�|e�24rz�+��v[q4�u��;���/fwC`W��:#v�=)XM;
OZ�ф�Mdp�Ez�8s�v/ �^\1�11���9�μS�*�j�=��P�h�ڰqc$��|�0a1Ǿu��l�]5U��W�N	UvΑ����t[��u,�[��݆X������
W�����BP���t�g���Q���������U㓖�55��[( ��'𛗺��+@ݷ�oxvC����[i�h��W���<��$�WFrRSS���)X��
q��f+#J�MG'`ƕܽy�Ъ}û|.Rn�����s�c	mL���O{遑���"%��Z�MNr��� U� �	1��P �]<��]{�:�U����5n��w1���/��}�3�N#(�����G)��E`���u4�쌠���#g+ƻ�M�6���6�~���/ U׹[-��Xa-�n��,p���q>��H�����p���n���|�흵�#y�I5���=H`�烶i�x"Vz�{���*��5��,��^+�0^���x#���GRK< �K�H=��0}�`��M χ�T1�,pn�6�ɇ}�U0 �,�*��r�i��7��'���O;��"����:SD�#o�N���?�k�=�NEacv�I�V(��i���Կy�rL)ҮP�iP�����,�95��3�
����j�2��OH��Q���ps��ߜk����5R+.�&f�o�q1x��O�a�������uX֟�Ь9nv�9̩��`���g��>�3*����U0@���5�'�).O��V�����K��Y
=�d� lp�o6�c ���1(�yu�j�-�_`�|"���׏��ju/������P�jDh���r1L_ۨh:�v4��"��o��3����i2
����ZV���Iؓ��	������L4����!�F`���Pa�"`��@����Eaq��*���0��t�08�{T[�2����7�Y��hh����P׳��^�>��p]��O��6I���З������������ORR  <���x�6�]�/�֩M=)1l|q�AV�B�x�`GMgR�˳(��㛟��N����V�.�/|P`r�,Z�򌊒����?E
i�eVQ�� iD�R��7��U�����c޴�ǒ��_{�3_�$4�M�]Pq�藋�����'X.��l.�`�տ��=l�5!N��2���^Q7�F|��+V�z�� %��$��q�����3z�9_��%�)ť��a�7P�������������O����M�*��e�j顱�����ر�<S���4��Q$�֟�>�̖r��%��A� 5���?��r�Tc4�՘:����B�=��Ӕ�	c�C���}�(�K��a���;���m݃�1�6f�'�������sS=6�B9��Wd�+C|�!  �\n�um`���QJ0Kg�)����u�?��`Z�'զA������DK���֖��;��]����þ�7ﴚ������0m�����b9���(�jĸ�f����[>z�+�7�5w�D�r���L�
'?H��4u��*�m��-��d�d�q�oo�\\�"�Z��n.n���u��\�����%�_��md��H�zθb���^C\ؚ!`(3@����6��/�XT���ݶ�8-\��AXr����)��+]�����bϵ���3�
);�*v��n���Ou��I�T�K����'q*����)o�[h���E������h������N�{�������I"-}\�ϴ߻�x�/��ل�#�]��/�s��\~���H�ԗsw�$�.-��h3e���9�.��8���3��o}�}W�ǜ����+o����I]��HUV�c9"$9����C��+�� ����
�̢1>�Bݰ��d>��ޙ u����3����*��
B���=����r#D�T�j:��3������*��H�B��V�p����.�8�����ֲC��ˁ���*!��:�YG�(����s��J��h��K��9k0��_Ph�~h�,ޟ�:��
3�0+%�u���?�`ʶ{��I�V�<��֑$3\���j8�t���m0'�G��kY�!z_K+�G�NDa�N����4��`^�%�>V�r[i�r��7���i��yy��If�p�i@x-��ל�O�a����Ik���ϥ�<��,%y�or)]}���__c�+?t�����Z�qc�&�93V�r\�0(:�5��Wz37[e��-�N/��=2.�����Â��}7F0���-�+;�����jp����~�0?�=7�G�%��0��s9��Wp�6Y⟅��;p��n)��#�==hɭ2��ΟV��T*�5�`�� ��O�ֳ�ʔݗ�̔@�K�����ۼ4�l�s��|&�IXE���8�4X�~���ۃ�j�G���O�O��&��H�ܨH��L�kC4d�/�g��~¡�?)R
�rf���?D� w�2V��[4��R<�����2�����0{��6����f'�8R5��\	�/Oh[��rD�E!}���날0:�a��]O�W���7}���v� ʎ[�o��n��[���yW��yL�Q`��
�����s���6�8��*�y�F��
��ǡ�yx����H6ޣ��M8��J��`5�r�5j�a�.!!�ӒX8�<��DI�wI/(�s2	�ș�;r�����P��	fɌ�����{wK}m�����Hf����%�&/:��F����.�JQ�.�߶.���xm�[���U�%���G�{���b�fC�%�3cG�.J�U�m���F�8�Eݾ�c�W@��6=�5c�_��ud3���+8'�$�R��4׊�I%Nن?#ȸ�]�9Z�և��<3��k�����G��=Z�ų|��s52b�G���6K�(g5��KS&1ς\߫x|�ٽ�O[��kG]--�a���s¸t�v�oL���+�#���˭/�3�$!+4;�?�O%��ʹՑ4�@�U��߫���䴥!�P���{傣��0W�&�FE��{�+Q��<-��TӶf�	'D��vy����'ɒ��DhE	�x�r�sS8�&�p�IY��8<�E�}�.�����������^�f�h��< ��uҙTa������ 
�J�Z�ޮ����b[�JƎ�TD��_�J)3Y���.���6�~/ّ��n��B�.��߆���BKK)rM%�$N���&�:C����?���'?[\m?����0���Y��;4�6��˵6W�VŴW�{�s��r��۰�f�u�fʀ #��8�p���8v�+�ٛ�k)������~�2��?09a
X���Y�$��y�&Kʺa�V�����aB�k'�4���ҟX�&u*4��;9�z&!�$��%n�b�,��,�^�d����XN��Zxq�WeƧ���IH�7�IG�����F�K�����Z��V��F�]RsAc`�O`&F0f(���N;9x"������x���>*�e���O��{@F3�Xٍ�'�+�+��kކ�zї���r^H�3_8	<���ݥ����Y��{���)�G`U+�+y6�������uIj "3TL���=�\>*�PZ[m�\%�f��䲸@�k�?�Rµ��^�uf�����|-s&����c28���_Lr�W�������؍Z����U�Q��@�L���P��@T��;�ɺ��Nʳ�5L��h���%h�a|��D��8,P���q��0q����S2�vҌyZ�<ه�K\��_��3�I��D�o�>�`ܔ���#�S� ��R��]m
C��7�}0�ZzntS�@e�i�7šK4��.��◙w�Fy�{ͩ���/�Q\�����ℯ�Cр�A���O�
��3��dYouV%{��6�b
�ħ��=�XT�ֻsR)�[^�8i��į���P�%�W^�6�p����E���Z�m��nz=y��֋�,���P��!�UVQ���,���;<���w~,���&�n�}��[:�+	�Z��T:"���0����H�9�#'!L�g��Uy�:'^C{��*�{��dv�#2hu��ׇ}�I�Vx&���M����ށ4'��Bl�+��>�DG����"���<9�׆R�9�Y����%$vɧy��LW�Ԙ(�0ʯB��>C��rS�V�y���H�yz����m�	>sԹ�{v�@c��-� ~� !��qZ��ឬi�s��������dZW��:�ˀp���]!�o����XKG����zM��a{[�� B-�/YSAu�P.����-ﾸ}��@S�9]:;��[�Z��^�?=�[9Ғό���Yh�9��I}�/�`�)%�7CGK�Elg������8ΜtO�+�3�$=
�-LaՉ��ԍ�r
&)�C=Ce�(�g��X�Ĩ�#�JVb�1�9�G��t��

f���Z��U�Q�$�R�p���şh�.�� gk<��Q����*�:���gf�A�qVV����*����M��k�v溎���g��[�<d�wSwN��R�u=27�&��Q�؁���Ղ2�&r2
�I�q`6o"��-�#&�+S�*��&��"�������j�����|aQ�^��Ke"N�Q���WH(�.���(Ֆ\M�G}ڠ(:Yf������9��۔�wZ��˅v_�1��G���|��	�[�h)Ci�'+t����կ�N87{�����HKP�)�^�bFU%�����ɕ���d�Q$-.K��8+�#�v�6//��*��2�-ζ����ssO����L��9/(��O�P��e���T��q��(�0�,�`ʫ���A�E�ן1h��ge��I����>Y�w��^b�W�f i���ӭ/=��T٘5�e�l���)KƔ���@�m���5�z�ZD�:�җ��|�Wc?���k�L\��v��\���?zu
?��wF[�yG�֟�	�����Rº_�$lF���5�����;���Il�7}���~��m��9�o�bD�����(����7�&��F�A�����qp��'=�d��/%�Ȣ]m�F �G�wG5,oGQ�!*"�{��i�A�Z���T�H�ޥw�.-��	:�@B��z�����ywfg�gvvv���)��4���#/T?��YP?D�܇'܇�W�)���O3�;��\�j�Eji0��c�(ƽ����E�G����8�8sD��kܝ
�w�x�z�����F��{p�'K�Ҩ�㒴���
E�����q���3I�P3l�}h����R:����yVN\����ٖ]�7򧔜��:�Ѕ�������cM�Ie��5Q�k'��"j'�Is�a��煗!��nV���I�e+}˜��>/�fO?��}C�$����K���*�?
j�p���rY�I��{�Lȱ�\k��@n�f�Tm%W���ǳ�T�)�% [s�#ۋ��-BF���y�'Di��T/����m���WV�g�?p�C�]t{_�y��7K$���
��cb�t��p�ְ{�w�����))��d��g�>�o-
�g�J=�z4*o���5ո8��j�H!m9�#���&��z�).������xJ~]� <�ĬC���B��P����U�`<|��)j�we&��UI5�a�{���Σ���f�>�M��w��|��w�l8$i�
��� ʨ�A|�� ��X�[��z�?�76c����V���.J��y���ā@`_����l&��ܜj]���CU�_:)灱<�����,�;��'����''���e�����)ۀђE�)^J�4��i3.�&�Tx������p��^(�Y����[�/�
`뚷��5�6�L��I���zF+�㮍�8���aIj�$V�bb�x������m?��ST�U�ح�)hv-�b���r@$K��K�4ur�&C��F*�yvX&Y3�j�FuI�����]�{}�粙��Gռ4������߈��w���]�ﾨW!���~C�婟�'�:5��}q���r�Y�`�����ƲJ�E^����aB�>�8��܍%<5�K�H��vSf�P�rq�����q���%.y�l~N�l�$Ӄۚ\.����+ȣ�wۗ<��q������#:�uΊ`z/�y�\]ui�%[��ϱF�27�q���r�(m[?�^��k�GU�<��b�sdEݏ�2�&Ҕ�o�%��~PQ�H_R�Ux:`5��A�奘������3j�ۋ���25�cc�M}�J7��^�5�0}� _[���K.�ރ*	��0?z�l��䤞�0�K�'�{3�P���?�����0�i����]}�&�B�+�	&��5��n\�/�)�m��&RFiT��n d�F�ce�ԏ
.��[\�0��Mc�v�l�(����f#���a1����1�
W�v�ZY�F§���i�\��s �������03�M�'1��uf/����Uji�[������5���6L�¼�ST�m'/d�}�����{��wĿ|��'���@5���+�b<�J��mF���m�Q�}�	�Q3���2�d_��18��0�Al��$�z1eĉ(��R+��B�A���.�Wy:ځ6��?quƓ}w�A�e}�Y�)��]�O�İW�S�=V�'B��F�d�at^6��l�{�o+�w?�Y����y����>���cͤ�Ev:6����>�����(u�2\0�O>B���D�^
� ���6Afc=�K�폸D�y��?��;E+ʇ�=8Ӓ��R;���V:�⺴}�_,Z���6c�� D��fK�ɱ>�����{S3�6�"0̋�i�U7�wu��[��r���MDQ�_��a^6�o=͐��c�S�{k9��e���&T��e��>�J�Y������zñ�~�K[v>Znt{�s�g��^rޏ��~��:�֧�ێMv��k	]j{����G[]-��[x�K�A|(]�Կ_�c�Ks����Pţrw�#8tw;����<'�J�T6��U��~�Q-黁���D�R��hco�:���q9�_ ��]w��V����wZ�4$ �vzf!_�����7�h���Gik�t �AEW_����tY[Vd�����Dn7���pp�M`~E��n�O�,'��#{,_On0�u{`�ǈټ�󩔟�Gʵ�v���
��8��~،��:�����\�fk��j�#NU$*�|O=��b����'��J��9מTS~@�]�����:O�4�ɴ���v���M�g�mi�̛�F�Yٙ�Q��O����\�`%-Q2�pG�������ff�t�(*�ғb��	�Uĩ7,U�y�2���gI��4�K�$�{��ߒ��_x�pZ����B�D�v��a�
�V�5�~Â�&p���qj���W�;5mJ��;��.�S���>FO��d�Sֺ��r?c��գn(+ۉ��0,}��@�bZ�<^`�J��d��f�壎q�� Y 6Vx�Jᓐmi�+�&i�w��t����j#�J4�WzȊ[��zwF���R#�d�,ҧ۪�����%D^�K�� �cU^��`���@|<s%ӵ��Y*�����MU�WuXQZ���y'�S��t�z��$� S���{��Sw
��F߆J4�P�6�-HY�k �1�J�/.-��~4v��7r�K�]������1Cnh�Ä��䤈,D���r{ES\��p\]��XW������Oa�vR�`�~��C�;��>c�'HN�ʉ�G�p����O	Xa?��x��Wm��l����M9� f��n��q������c੻N��GH(��m�|-p$HQ'j%��s�R�#]~p$x�i1~F�v��J�J�u�ޣ�ʛ���b�[��'���M�Q�	���h�xz� $Q�h�`tZ���k!�O�F�c��Im=�S,�`�����;e\C����]H�'EWP�o,̜z8{=��Q<X�ص;�z����B�>_o���tI�g�6�S�/t��ɴ,m��DPB�����0�ǌ�M�T�,<be���'�C�<�Z"�]8����E��wJ9�L
���z���Y�B��e����
k�s�H���-�kዙ�o6'�U��'��J���Y�#��d�bz��j�9o�.���|���H�E�ӝ���x"���
����UڿJ��_��W7�����'��w�,Ʃ�md���� {J�V��y��o��]n�r�"I)�ߛ�`��� �ɴ��w��
[0�ri>N���k.�u~��m�]7������S�V+�29��N0ǹ]*̬}_��7*ot��]�="���J6���K�WC4�e;����s�GFlnZ�y��پ�󝡮�n�b�\���+�=MK i3:�v�����~�Ej�:a���ꐫ�x�;<���ߴ��:E=S�r�ޫ�ې�;��Ϲ8� �(���F���x.�n�א@	���ﱰo���x���:fA�iԼ��x�"Nx�gK�7�É+��A���F���V���&�V�M�����6p�US��G�2���<^L�Ok���Ѫ
�\Vr���f���0菸�2Tb#ۆuq�c,<�Ⅸx�����l�.̱12�DwU���220��Ot�9���G/H~5v�uҦC7U�_�[-����M��-��yĚ{��eD�lu�zoEj	a���Z?�k�ۨQY~sn|e�,�(U,��CL���YJ���@��=	�e4V�h��vJ�,��-�� �G�Q+�
x&��K%\��5������P�/���X���g�����W�,*0�H����-�}軑����t����M��|yI#�B�Z�����'�;���8�Z�y*�n �H�*���P%=o5�gl$��ߩy��=�%�T����L2$�zq08J�"��{�;��pmtl�z�vl|���N�B$5�����U@����b)��k�Z��
�	:-'�Ń�ӣ����ǭ��ʣ���]"g�J�6�LE�jؗ�z��P��6�S��4�'�ږ�.�8�ԢE�oE�c��A�ߣ=�!�,�E05HT>��-��-1�D��V�8��Ʋ�O�#vA�-��|��FJ,�?e}{,8���92�zAd}y�k+K��W�o�<-��.�K�U����|?�`��y�~b��jgL��A#$�Fq��^ad���5����*��������^Qc��HIDp'p7���BQ��A�[g�C�{r�^�Gc�M���2��E�nyO��LN���~����B �����20cn���k���-벗�~O���k]68��~��T���"���-I�u���,,@J�G�`���<�~�i����:̱>7�]C�t������qY@%����m��a�:�� *�?f�oC"\�=���*D�ۗn*U\�7��G�	�"�o�/����X�Cv<� yF�\�s1�[���V��Z��O�c��fȝ�B<ju?`��L�Qry���R���y[u��n������m},���<(!�� X����ܕ� �U}�}���8z3��4_F_�?��~���K���g��d�=K��U1G^�� ,S��[/�"ڻ��K �
��&��_3}��/&���v�
i��iK�����ۏ�G��G��2�B4(����t'yy���bkř/�.���D��:���z#(��h>��V\2��j�jO�� q2�L��ωg�ضPѣ���>�-�x��pz��к_Ǖ$����u�	��"r�t���~�����4\}j�q�{�����k�Δ��XKy�CyQ��6f�t�nM�&dhh�������D�W�k�~�fY�l�;�a�0��8���Ɵn&%�8�NM��'<P_}v�?s���8��J����t6h�:�YY�	�o�G&pCȶ*���=���s��J2�z�|��θ��!Y$)��	.n�Y��8 �9x�/�	,���{m��2�k..;�O���H�����S	;)�DTz/��F��b��J�N�t�RW��2�㣗-�K�,��d8��T�Ƹ	����F��S���p��IY
���X�(tw��17����wf�W�83����҄N�{P�㎉K��+ױk|��Q���߱<@J���9J������,՛cn66jRm@$ ����5�)���E�d�~�jdQ��Aȇ(X����ht:����ΟV��*u��Xw+���n�/m��*�I������S�*	�Q���A�o���a�o�^|Ϧ����M=�t�������zuD��Q�X��K������eߊ�4��_ؔ��5�4���,�=ٴW,��k��h� ���<�����/O��G�>
e��;΅�����JW��;Fy���m�(�!���p�`�X^gae�L�Jf?ft��]�<�k�UꐚyՐ{z�0�f߸��2��:�8�B�jB��y\�#�? ��	򂥂�*a5�0��1��W���(~p|9���&�Γ���ԋ�4�5r��óhC�؍��|���Y�V�^��^b�]�q�l1�d"\�d:��P��Z�tO@Vc��+̷皅rH�P��J�nw���X,G��bf7�<Fp
<߄�^��d#D��=�+Ƅ�Nd��t�`�mr�th�/|��H����@\U>'{d�BF*fy��^�MH���2�2.pB�ۨhP�	2Y]]ujrFV�&u�;�������_�!�ˠ5Xi!N�������T�C;��o�ު���?�+�t"�"�Ht7����!Ԏ�}��t�{\�������H��ў~(z*�'�#����G���µ�{��r]�-���c�L���2�%MB<����:�A�Ҹ�9U���C��Ћ�D��X�_՚`s?����4�����;�sY	�0ϩ.V�/�f�#X�Ao� O�Z&�9�jt�e.h��OD���}p��qaA�rC5��ZP���u^�*3��;9EE����������f����I�&DW�>Ey��Wz�uK��x���Q�Q "�s��Զ�4�q؇cG��L#g%�$�+I�B7Mٷ��2抴�������cS����?�#�������N�n�Z	d��/Flj%@�Jǒ>Uѭd��@S��4�����m�U^�f����Ǭ>���AN-Z'�38�)�c{����	K�'+���)���/�U�3���ӄ�߀O{F��:��[E֚ф~],,�:U:��y�a�R��ԋ��.ʧ�V�0��DK0K�%)D<n�x�I�`�T��Q�Z8K��l�d�Ȭ��i*���7EA��� �;P�qS�M�D&5��U=�W)�$��1���>/��t]��+�#���Wu�nRN�X]-������ʟ��8X���X��(��|�[��4��̪���;�񱁡��GL����s�{є9�����"]��. ���w�(�\P�%<M>���GtG�L����cR�L?]��MM��h ?˽m������t��j��/�P�B̋G�xN�n��x�
xF� �L���D{��������~�!�
�X���߶����q���>����sӕ����qF�B�J�u���O��1���9h���>����
��������1�Wl	���&�%�-�?�5k�y�8�E����YŃ���J�ҿ�H_�!���"����	S�Z�Udt�|��h[C���`���xw�����	dS��V��}���Q�=���@]@ʗ
��{��`�?G
(��`	#�ٻ����C���R�h����,���
�4� G꧞rf
�L�� �#�8�7m;�p�#x�u�f�����*���]+y�s����cI�d�<F�O=�F����ؙO3�$ć�X�׭��+,����;ի8..���M�R�����z�J�Y9H�kJ�����e[��!�����{N'��-�]R���L�/�3M�݇s�v�_��l�g�[�~ֱ�>N'��Qت�����aS˙�����<����_��9j@�\%�v�����ڍZ���O�+<�ce�n�?V�Rcd0Z�t$��z#?�Ć���	#�ء�E���1�,��XM����|�0�����1)j��ZcaqzP�������Wn��C�<v�2��+)�7)�=���Q�xk4h��SK[�AU��j�b����|t:*��-3K��Bf�c��	0����{���5�/�nA͛/�����>��Ջ�`���0�~�*ӵ")�-�X���~���}�W/��0Y��c��e
�!l�l����Rk��h}�ξ�����ĳ��1""��^Q�U���ߠ���=� ����f�<taE@%��H������B������p�8���3��F�B�bAmՙ4�SZ���ud�y����$�͌'O33�j�Zeq2����4~Tq��u�G�4c��]l��M��!�}O�a��x��+��	�d]�;��rz/M!�Z��nj1]ǺΧ��ΩqG` jkp`ղ��EUj���/%� ���\��S�us�IL�n7� ԠN�L^>f-2nzy���tR����|�:Ǵq2qK7�����#���/_���|�6;����q<V����i����{.pȨT�k�>�`�_S?��|zz��(�N]I��c{��-�0恺:Y�S��:�,���\"� ��;,?����	�2g��si���,2�_�c��lm�ݘ�W�N��٥g��X[�B۲��O���;�	A(��veNk�aDW۽����V�85�y'r����t��Q�Dۡ��㨬�����9A�r�R��]Y!���=B6�k�H�i����`~�-q��s&�@��Ε��-(ؼ5,>_I��2��x�Ѹ�1���#���g$��K�Iڈ
���sE���3��6���g��z��xa[u��[}�B�,A�v��w�_��{��S�Jk�e<�������P8p�*Oe�v*MM�95����h�Ё�m��YT�x<�'hy2=����u�y^9�Lw��I
�9E�r���;�[O��:�TU�::�u�l����[��* ܕ�I����9YO�����o�s~��C���>�5�[�r��T���2�U#�#��{��8�J����2陙�F	ɛIA�RI��C��&�t�h7n��`ƚU��{�d<��i*����=�{��wre���x�����������d�
"�5��.k���o�Y��TMڣT��3
 �����.e��������BBd,�o��H
C*՛�9^�2���-����(�#zG����Bj��n#����ÛJbm=t�9Uboj���v��r�mtn�n��h��I�x�X���\ZE1�_��W�����1L��Պ͎=������*��Rg=`����(�4(�b�/b����<�n����ߵ9�1�����J��AYV֌��m6�R�O ��n�Jh%p)��Cq�����9�<NXg.�S���%�l�� 	g�|���!t�+�G���U�ǘ������o���cP��sԖ�t�7����?1��Lͯ/���xmf�eE|K�MH����M�Eu�1�������������s�7:�y�&z+��	���&�)I �a�e3��M��N��	�G�����yh��I-���n�)_^�.��_�N�HU�2Y=>�i�a]W��&���ӚX��C{�%ƙ���	6�Jes��!#���NEU��lA�J6n�gvM�5�1��E�M��,u��ӎ�G@��S��%���_�d�TR�=��a���?���ش�0T���Z]-���(JO%+��Sbd-�3�KV��f\\��ս]�-���5�)�g�k˺Uj-�$��P�����^RD^�� �Ewd�`�ը-b���\���K4mrˏ-�҄����Ϲ%���키��3inɑ�e��9�����z��S�f�U{euX%��H���zW�1w��`���T���#���2��L�x�X�m��'�Ib����u*�{���}s��������b�Pj�5!a�5��+e�#� ��'y��"�z�i=���r���8���
>��$$2���y�T��7�I!.Oj7�="�'��!�}�[�������CA������o�;A�x�8j^	�j�@��O�����7��d~�v���U7^.�)�oԲA9�'|�k7	Ս-���IIG�p|�틙�-t5��0�,�N�ڪI;>������`�7o�����C�yས*����5?���ϡp�>y�����n�xJ��J�9L�9a���Y�q#���m�d�FsT017#ci�X5��GCR����ҵ�KX�,�/�c(ҳ�p�El�+����Uo�ya1�"�N��������XA?�Tt�M���1Ln�Ś���篨A�:�е㙄<䗛�I��,��>���x��9=}�gm��ǁ �n8��.OLZ�b�BQy�	�=yvL��>g����乹o�	��d-�>j�+��٫������S\��d�����S=��Ft��gϊ}%ΐ�Bl�&_��B��3�me��DnI��Ԗ���O&k�#3��N��L�����N���de���Q~[g)�Ȕ��NX�lZ�q��|�5��{��ߥ����X�a�4�& _�;���ݐV^���d��{~)a|��G{s���"��x2.�7"��8L���FH�AznC������C#q[2*B?���L�����tt�n�X����@�&n�#�)���g�C�e�WbB䐈B���v}���6�Q����^v�s��1�TR_L7N�U�����uzs.�����ߓ5Q>���}g�4}eKG;o���Y���;�[���2X��� _UJ�O�=�v��D���#+=Y�n�:܇�oXs�,�z�>$��/'����&�3�z�魕Z����"w�Ǿ\�'����|��C�ε&S8�kK�|<{�g�M󹘙�!F}b��֒�B6��?�.Ύ�K���Y�|��[b���z��¯���o�;dhsⓖ���.��v���;>�1A��N�ط~�6���||��z��B�ήF �uos��{�\A���U]'�!{K�g�o�����a�#em�37��������h�7��
�j�	��:
�l��#�Z\rl��3ض:�r����{���M�K��_��sRY����ϫ��� lGR9B�1-3C[�ESDY% �rG���#/���*��t.�:�&ZR��s�� �X[�쯌?o�I�J��\X-7��7�E^[G�?ܟxe�f�N"3a�1�mG�(UD_jF�Iߚk�t�}3+e�FnV����>m#^�)��g����d���O�@FJ�"����1�7f#i�A
e�Lӑ�Sb�o����:?.�ن��kt�7'�֊}�uB2u���o!FW�!2�(E]���޸��0CȮ��zX��G��Ҵ�=�Zl�N:��S��w�����M�2�"(���x��DL�%J�K3�;S�������:~g�j�Z(��%'C�[�l0Λ����	�����Ī���/��7Q�B��}�e�I���!�Nf�6Yg������wH͖k�s9>,}�F��r7jȽ9H����]VY���R~ਫ਼_�ŝ>O��5������~��Rwo��Q��U/�R��Y�H4}��5YW��ZXG����_�}���=8����Ibmy��9�}�3	m��� 5��B�4��Ņ�D�
�OV�����빆'����6�8�5)"N\{�l;�#�W����C�`!A��z+�I���=	��Ӏ�<�/���<E�����zI@��(%�qW�G9�^��G�����$�)(*f��uv�P��z��ǀ��:��T�Q���,i�Š��X]a�Jh���T���~pZ��C�|��L~�^Zl���$�J<<|O�2�y���~@�i�<o�b�����.�� b���V����g	�)��R\��R��?L����b����қ����g̍�Qe�
���z��������Ӈ�5��������cW�'��,E��H���a��x��������ꙅ���>�Bt(� b+�>��|�~�Ɗ�8L�-��� 7�7�Ρ�i�� Y[��[�%��Σ}0;�`�<?  �[i��׼%����ܱP�V�����4YL{�*t�B�:o�����
����_ދ42�����&��E����"Ջ;f3�����(}�BӔ�/��L�H�F^�ƕt�AN�!�ƨ�`���,�lu<���El�XuZ�[4�o}�I*��!�?�{-��)�B���q�Mt���&_<}A��� L;#�;r�����dB��,t��!#�#��0��yxx>���NV,�C(���Q�`�"i��UO��Yƕ56�wF�f��LҨ�[Y�1?coB;1�\��,�[�y+`�}��qV+�4ASu�K�X�j,�}P7$�.��\�97�-.O���{�i�S&*��I�Q��̈́~65��`����NT뷛+��a������f����q�Av5����W��}�}Cvq�o��xg��-����;{z���bR��l���cR��Ú���d^3��J���$ZUѱC ,N��E�������b:�i����C%��m�<�Sp���٦(Og�l����5��V:d%Њ�0z+��9����� (�����Jc��9uXE�[Pa�i�(
)?��K��h*�D���g��q�\�6hT��J.u��F��7f\ʉo-5��짣����1�&z��B���5��Rꅝ�vV
G"MB�lo��ʮ��Xq�j�����z�,10�Ǎ�u��K�R�O���fy��2����t-����?�ƛ�6��i�O�B���+Y�ף���7ڠ�[�
�'w]��������W���������|�ÈE���*=O(zꃗ=�59�(M�̼o�A_�)1���Sl�t;s�(�:�Ąg{��nBH�YԖ�.�}���KN�Ly�>�!Eܘ����Fvca����7ak��(<�-�G����P�����UȎ��;{>�]?����Ԃ���� �����WZ��Q��%�
ܭ�k%ޝr�m�!�v���\�B�갳�����VH���6G���95&�÷�n}��U�=�?J3=hse���G_HCv��^ta�/�>da.�`<�]��[g�����<'����oY�b��&��c��q{�+/[��!���"�O�O�胄�	N����1�>m��^��7���OӢ�6*�eU��FC�|�٤d�0�@&(B@.ta��~��hn,��J�y6C�Eء%�A���~Z*�����./���H�a5��^U51�<��0(���L�: ���K�BV���٣����3�a�y�װ����e��3�
�?�k�o�twrY�w���.?Uf������-jHZ�xe���TNp��z�2^\:�F�'P�4V�=4Ō7'|�e��Źr�=�k�7��PX�~*���w�*��j:Ew"\<�\�j5u�a��Ԣ ��|��r?�8�yM�r�:A/����ϣ�ˆ9՛	�x�f���f+���4?�O�دE��=�U�aQh�\���yᐰ�=���]П�~1J{���5�����2L��M���*nB�� Xު�; ��'���϶;��n�g�}E"����${�%��q��m�<�r�j��A��ŝ=B��D�m�g�}�e��)��I<�ԆD�H�TE����i��gX����.��,��%\��[�y��#�>�x�#��?�L|�N�>�|�Q���Գ{��#��p�*RV	N3 ��V���3��&���^0T���>!k(Б_�����}��Zz76�,��l��#���7\��'yP���KH�p'H[��O�:vv��7;/�;��Ls:MNӮ��=����_���D�5bM(23৪�nʖk�ۢy���x �78I��G��=�^�O� ��5�>��?�����h~{��r�|q����գ�Ї�0Y���k���iX����;���/C[R,ʟ�������'w���o��b_n�*n�\)�d�UD����ԟ%��pulB2�"�o�m�BpHp[G�܆���I]TPs���+Q��/�C(�u�	�dp�<��Vkn����~�ߦ�>���tu��s|������n����9eXU��<C}Fy]����Mb�َ��p�psY�[J,1��YW������֣�wv�z��\�'|�ȋ�Z�ev�gbbV2OE�]�$Q�O����l�+0���׻��1V��eou������\z��"-�tj��j	�������׽�1лfiX���͟Zn���c��2��K�sZ�}'z��=�Ý_i%���c}��4�.+|�06�zf�j4��]����DE��Lw����5��?��>���Q��V?�c��]d|mis.����(�)�To�X���ɓ��s���`RIos�z��,;Hk�)[�0طZ�'�i�j`�=^���㩽I��^OlPr�B�����c��4��=u��;�U��G˂�Gc2��F
2tw�2{���̗8�n��͎;��<���2n�d���ړ~
i�-�S�O^k���5�0x:�3�H�
C�ގ�?_�M��3���:0U*9%Vڦ������^Ȱ��/1v�(Ϟ��|�
MuR��������epa�Ԭ,CS?&�I���kR�}�QO��tY����&Hq�G���� �'Bt��*p�{#���(S���*l=��X���%�ֽ�7��ӈA�;�H��O=�P�4^��,2��~]$Xu��:Q���L��&F�,���Y���I����C� �#����0u�Z���ަ��-W�g)������<6��ď����~��{z<:u��5���~��"��)E6�>դ� /�,R���־Ar�C���Q�<��gj��h�P����iA$�4��(�y�S��*�V������z�?g�-'͗��P�%���+;ru�P�x͊]	���\�E��� �O��K5��_�;k��iy4�b��s�_D�ّ�~6
eK��9�9I;->�-���L���z.q,�:5��I�@ ��b�7gS�˼���vȮ��j���?�|��!Ӵ��޿�Z�3���ݫ�~��[ج�6�
H>���5ND��z�f<����N%g�FT+y����5u9{��yI��p��rS+���,7�6��1����~q�H����,?#<������|�Y���z�R�p�LI�d�BP�������D_Z���P�n�z�qv������y~v�ӑ2�y�H+Ɲ��}�V���0��u��$�ux�d�:G�֐�Ɠ~���<LNUai!�l�`p#ƫ��� �Z���p0�y	���g͗���(_3<>���cW�zJ-�I���3���4���*a}��삧�����Q���-�PJ��l�X80w����x���y��VR�x](/�"��/#�>�݊I-�o�e:K�q�xYz��#Lv��/�Y|���.��a��̍�͎�
<�0s�{� �o=���>H� �z�Z��ӕN�x����
�5Zi#`�톷Y��߉r�jo"q|Sz�����?�q�g��,��a�u�_�,�_m�/Lߛ(�����ȳr~�쾫�j�x�׍��fc�E�
!v�y:t���> $ţC���'��8t��T���c��1�{xo��<o������:���
H�3H�.�,����,O�+�/	)Ӽ�)z�n�HGo}�b������.'��Z�p8T���˨0�me�FYnT��bi|8��C09����.�(�[��g_&?��Z����k��eU�~)���Pb��* ����.�C4������g�pB�2aĜ�����T2��޴]���*/4Bc���s��`��T�X�T%�����B8�q��$'����Z,�a+���r�(m�[Sl(-�28ǉ{�L�=Տ�����u�?�������v���t ��汛�M���3�j��wb�l�uhk�����MT]��������h� �ܠ��5�|}�o�p���r��I��K���vH�,CC)2�����J�V&���~����ڡ��K �
.�N@߈B��ĕ�K��7���e�A�"�T�r?�?�M�㮃3FR(.f�mΖ���m��N�55����W����^Y_eZg���yI�]���-���P�Y��:�o�|Y��Eg&e��|9��}.�-����Q���u�	q۪L�)e�q\y��/^�%<��U7'�����E���R�*)�����2�E��u}뺁��{o@Ʀ�.RAm \(���♗���PH�=�@���S�s�A>�i�l�vF��83@�R�ߦ�ʯq���p��y�M{�ަ����^u�hԁ�9te���'3��4J�.C���405��iu�I�g���"R{orL%���xrϚ�؀�Q��׵c��k�_���ř�ea^�}l�'�QW6~9�}�ء��}��`�T���H0`�%EO���hj��=T�m��-��\B�M���ĺ넄^-+ݳZc�|=��72`D�?R$=�8�w���oް�ӊ��^(�� ����A��������4�ƣKetn��[�fQ��)�X�,�UT0�t�po�n��f;A�D�7{ۃ���me�s~��b������^I:AC)��IH9	���`#A�ag|p�����K���2�4��t��u� �{�C��@���Ѐ�4�o��E^8Y�̸{7�Al��k<��ͺ����s�l��#��>L�=Cэ��c6"�&����qmȅ������4�u�����E��!�0]d9�J��#b��
��3k����0��^`����Ή7�
XƻLK��d����#��xN��y�T���~p���G3����SvN'D�=՘6Zr��u�h�1X�iz��7��=��H!�
dca�i�u��Bc;�qO|��B�ܼRl���8��iV�v��C����b
�s~���7�{�IW�H&����Ԁ����~:��䬿W����:l�֍)D�S3���1�-�?9�d�ne�`X		璘��P\y�R�,*)�w7|���W3�0/��Np���&�S����K�$���H/�.�<�-��!����ͱn5�e�|�"�y�����+����|>�?�t���.j�P^H9k����s�eH�O9.����#��DC*��m��ނZ�,3퍱��f|@('a(c-�?�j�L(=��i٪���1��}�d�t}��5��o2-.=��j+����,�,�+��(�w���6�DԮ���4cf,VP<���|����B_EU5m\����,w��vi"Q����ԫＢAe��5$e����=�b�O�u ���^l_W�Q�mG�K R
��A~�R(~B�뻎�C��
,@�ʄ�i��-��0��~����{
D(J�ж�������a��b#O$ͧ�_OU࣭d�=&�1׼�ʘ)������{{[���W*��怷��,�b;�į��W�e�l�[Ԗ(��e�)�^����;����dl�=��q�LM='���(�^��d�qC��gO_�i���}/�l�(pD�Q��r;b\����&-��2�>���{c��IX�'u+��Wj���MtbR�����Q(������=��}C�"����Ե5��
�4�S#Xxk�Gգ�e�b��\��b��OJ�R���dzGػ����g��=���k��z����Mua:T�*�u����|ã
� U��,��Nj���� �|l7������4�x��e����VW��t�3S���2���Kd������Osz�O�Y�Ji�Blr2�͆���S����� �>z(�?�LF��5[� ״z>vt[�O7��C,�`�,	[����1�픥�ȱE]� h�>�<�7VK�6h�R��.��k%�<��&�)�ʟ�R^�Bk?�?���zU&̽;�hS%�3^���>�>_-7�c�o����>� ��M���YJ�RS'P�\�C�Y��Rq�FY)[b©H�ݿu��d�sY���J��l�f��2io�GH_y����f�>9J����oY����*Ý�����W��o�=��t�.o�G�8L�A�<$�"�R�3D���%6<ѵ�/Z�v��i�-Z�y��u�l
���)>���U�u��'�>��ʒ�Q�.{��"���|�p�լm�&�����IRɘ��X_����?����mk;�P�Q�RE�T�J	ET@@J�齆�G@zG�@h��;E�54��!�� ������d����}�^{�g=��M����?)��[��rA������a���BY��C.��٥�z���n�9|�%}���]�<�������1��"	�e��Cvvd.��*��V�A�V�j
�۬�UX5�X��A�Z��J�t8�ao�c�ĭ�ٍ}��,.�+Ysߖ������Q��J��H�}rȳ�<<|ښ���H^ �����>0��{R�,��5�̟6�n�iJ�NCW���?��y�!E�K�ͤ�M��ew�m����ţ�k�A/wTW9I�n���ez���褎���Ko!�=[7٭ln
��(��̌འ	���vM�B�	)��dd�{�<�5�	�&�Y�%;ߝݯ��pI��x3vކ`��D;�\0D>G@�{:J���[����kq9�<���o�IG�q����$��v8p{������s��C���ř�e�1e}��c0B��#\��9�C��x���6��V�����ԑvݜf�f�:`�G��	ܨ�-V�8 �!-��:=8�,�iS��,f�͟C��|?T?�Qz�����W?��k|�]E�����}�y�C�r�tX?��zN����=�,4n�0h�$�Q6�m�
����-�dŹtt�$7}�����E�K4Y����²�Q�w��I9���?�����2��s!ڙ��2�����d���8F�� ���͐����"�(��f�,#��+)�o�3��r��A�=�$3�(�D
[��Ӹ&B��%c:|3�+�N�54Iı5�F��\�aDD>�5�.�m�Z1����׽h�?��^��P �!&<z0�#��k�d]һ�pl�=�V�i���Yi�ɸ��ﶚ��u��hLM��񖍑�_�5��(�O��q�ʬ3��/�kɆy��#��ڗ��+��sp�T�SX��b�%S���jF�֜gd��}~�%g1����O��~7����m�[!�8��]r���e���~��W
���$�wonҧ�$ҽ����m�YS$�X����n{���Z���[sΡ�G}����/�g�\Y��^��j"HX�a��2ν��@�"+��$�X��s�)d�O*`�����f]=A�Â���� /ҫ�d��_\��gGt)ș�;P"�(��~�>���tYxI����ki.����*k�_n�'�H��Bf�i��*���%l�����r[�1��m���I��_/tϯ�J���.}�s��ю})�G�ܽe�4�M�����Yo0��yi%_����uV�a1���%�R�ğd��W�s�_����׳���$ٴ��w}�����.��rf���aH�Q�$���yh+�Q꥿�t������J��� ���^�"�x��?��F��5���"�G�޸�yt;nG)�\�+S��8g�÷�f�z�M ֻA��q���3/�%E�[?o�7խJ��w'd	{�>�btz�dE|Ԙ����_^4�	���ݖ|%��C�����锫���ۙ������I��-P��%,L�� _E�Ωoz�8%�.;A���G^���I��8�O��Yr~���m����QV�R���\��P�m�#�a��XP ���.�0�N�-���U�������  ί�<
�=t�F��K2�4��ˁ�!�>!�6�*��(� �k�V�8�;���߆�7��J��~ћ*w*}ǊE��i�˼�Ţ�Z�t,�]m5��8��Z�yנ�-��1Dk>���t~��8}$�Z&&������ z/����("��G��=����q�6���f��tE.D�$��K�Х��j���I��������5��"��$Ʌ���J;�Q��<����c\ύ�5�+�#-�9qRFfC���?敕�n���y.rd�wo�z�IIAy�]V<�bL,{/:��&6�����6r���2�~C�E< !2#h���r$��"Zr	b�Ks^���(���ة�u~�nx��FI��O� ��oGG��$���vr_P'��1����-kQ�#�ǲ�u����w����Z�K�����o� Jϻ+�1�3*NNk�m%�oi��2nH�_l�bİ�o/�M��X+�Pߴ;��@2��z���T�~�����NZѣ��cV�ߕ�^'�I��/S,&�G�[@��\Rd���s`_(�s4�o��|�.�Dz:�z��@{=q��.~��pn�*@�E���t/�y#[y���1nN�l�.=Zػ��Ѣi $�:���^�����z�r�AC���Ĳ���H�~O�҅iJ�j�fT�S)㥴�RHW�v>6�brz�q*Y#;X�`���]��"�$�d)��1Y�O/����j��C�tKoIlq �?��G ��eD<�n�1�Q�-՞��f�9���$h��8	��(s^s�u�ۇ�����m07�T��I��-���eXPlo��R�~9���%J�^���4�B��4w<��&���ʥ��O���&0P*��[�N�R��$�bM��t�p�vq�L4>Q��W�h#$7b�%��)�?����G���(R-�a��4AdI0�O�j�i�"8�]��������X$8h^=��Cnl(��QE�P'x#<jL5M��W�n��4Nk+L㝔N�g�ǮȾ}^����t�D8�X���K�57Y��A�y"V�1n�o���B)j=��!S�g�5�S�f���B�(Q�U|6�9Y>��W��
�HΗ�i�M�N�ITGE�F@O?v2+��t~E�� j޻�c;,Q���}�P�Oh�$ev� G�Qؿ�صI�]|lt
�4��.PƷ�:4d=�=q�����"yT�ҫ��z�LT�� �w����	q���/������{�F�n{�nմ3�dij�J���3����Q,H�^jYʠU�+��x�(T@ܕn���:���4}d��h�r���i����M�ĬD:h��2����M_0yO�!N�h
�V �צSߏ0�_��sE8 -�=c�Ԥ!ą0!Lo��xi}�n���4�m��9�G��k~�O�G�w�r3-�ɥ6�wڨ	�z�yn��L�_�T����W��u���V�0�K��xN�6	�
�+������sHFm��3�D�O���}&�9�i������ߖ6	PyL^�@J���=��N#Q�oG�O'+���x�I�A<��LB[��������'��*�������9X%^i�ihR[B�[��9E5/�z$/m�,{����6�	��p�`e$�/(В�=��&����J�ҫ����`�m�FŹ;�M���i�5�C��,Ύ���p=�����I-���9� w�"���fg♡�K�͟%��K�Op(��H�v�bHd���A����u_ӽ��������J��נ�k��,���#��W��M��z�nh�reE�0b���j����	��I��|�g�B��i��P#�x�ō!�������� AaꃄG�dWW+�������u�[a.��b�R���������EXM�4_ƭ)���p�X��3i��� ��ul�<1| �aIA��� �����"�x�4��{�C4�採�,��鎪V
����+Ŭ�F��,���z��ו��<�1��5�&7u��ARLoN��dվ�
}���Y�Z��hm_��rk[��i�kF҄���K�S��:����R����3�u��J--�-����
fb61�C����î�^#!���e�������|C����=���I�H��H�6«ղ���Q:�+�Rs�����&]��5��j�T�"�޽e���LU�}�����M��d?D^3	zf�|��fAP5i�Rg���/$
��<]��M0�f�������s7���g|���^\��!��-���F�������w3y�?�$if�7N�����K�P ]�2��~����Ʌ_R�U7��~BJ2)���ړs7>�� ͘WKal���m� �����OV�&��[Q��U�����\�6�h��7W6��	K�D�>��9�)��u��o�
[JJ���~⎾��*��e�8��+^[kS@*�����v���e齷Y�f�O�l��':���Q�S('k��n�X�n������2�v��]�rE����P��7��c���[�-���њ��Y�������GҤm�^J� ���'��I���zڽ�٬��黚9j߇����u�t< jڞ��%��C�}�Lr�#�r��H{YG8 ��J��7<�O%�ݎL{�>d���`M�q�o�GQ��g�6��T�9�Z�#���uqK�����*.�\����YU�������Q����tI>�r4�2�U�@�� /�i��|�E����V�K^K���oiJ3�IGE�=�`T�w����C���7m	�a�U����R���(�0����zV>~3�c��Hy�-�Zϋ&�o�D��#�.�RmM=�&�pP����i�n4���U���`c����Fq��������ĠL常�T1�:WH���i=O�B4��vU��8d���G�y�4YӶ�����hA���q�[�F"��D<�d�D7rҼs�?F���*a|�#�W����B�4�G��N�ɤN�ۙ3���W
ӯ����EH��le��3����ma�l������尼�����p�jAM��T���V��?cي���,��j\��a9��R������bS���>/��L��2.|�=	*�f���~���\��g�WH�/!�O��z�C3�Mw5�_U�)�����k�qz�� �w�(�2:۟�!yK���:u'�DWQrШ�m a����p�Ɋ�à8)�!m�%�}MpYɚ5|�CBH�P��4;�'s�'~�&�����M1�Ywp=I�saM��;�LBY�O,�OJY&z5�fq;�=�Y8O'����}�#mfXծ2�6L�䙛�k���;ه���C�#���r�F�W�~�R�L*&��-cu����^�ENJ���+�Vf�01��GS���sK�ŀv�5ި��Jo�OB��gz�m@��sR�R�a�o�⮉���������V�,լ�$�6o���)�3Q�U]mL~|�����E�5�W�[B��P��/�=���#������}��T<� ��g�x9` �1z�{Z/w}-�{O�GC0�g�
A8cڀ����[��P}�ej�2�r8�zt6�oD@�(��Ю1���9�����*�Ć��t�⃐�Y�-�dq6��N�"V����>]�;�ژGp��m�?��w����њQ�y^��bu���t�&Z^!�i"pP��l��F��'�(��I�=�p���=YWn;O!x2ڿ�j�Ϡ%���\H�a+xhl� ��v�Hװ`v��yekG���X���	|G�� {gXW�[`ʪPKNU�����9���"m�&����iճR�ס^��2��6m��I�e��OU���.��ZԶ->�t�,]'y�.M<t�~���	��}ż4��{��2(�[{2��to���颹��Ύ	K�_��I�ԫ~�:J>z�u�i�R��QŎqmh@"��m���J}$��q}(~��e9�{��v�Q �h��c������t��e�Nܳ�����ͤ� 1	w9.e�:�w�J�������fu?����,����֗aG�Bl\�� V痰�sF)���<�>�{��6�Tj�im�s=���C�6��X��AaATgTj$���7*m� �ֲe��9K���Ӛ	"%�jwa�B�PV{���fe Mm���+cw,%׹UvQ����R_2:�ʢ��[�t�?Q7z.�?�h�;&%�p��qّ>蹊���� �d�����Ɛ(�ٝN���K�t`��ߵ)��7���S���w謁-�8��mT�k����Ծ,AJ���{�T>�r�='������ص%�2C�<)�ʢ��5�
���=�Ho���@��Ź^��M�B)ߤ�̯��#�U��㕜z:��K˴�^��c��iO;%���T��7����r+ӌ�#�)��SE�^]�çP~��l����	�J&V#���6�� ���*+X�����Ķ��2@��=gi�s|��0暜�4ĩ�H2����a�;p�c�`m<���Y�W*�L��p6`8|��!�Ɓ7k%-��fvC_�����8��O��/�E�z�����d��jR�F�����z�[P�O�7�<�\#�N�~=;��o���0f��,i��Ke�^� \�ymO�3~p�H9�+@��9���+�%���(�i<��g4�=#��D�ē����ޡ���)?��뗾d��U3���M��]���y7���v�����-���;���ڵI"��]�i��u g;�S�����IO�f��u�m���Y����Xݽ��4�c�����O|M&�b{�	㥗V6�|Ps+n�S�𵌽$O'�8�%=���/���$6��Δ\�f��p�7�u�z-��յ�r���Ǖ��y_޺�	,*�(��B�1�n���3��o����ǓuN�{6
��vu#�i�����7���?kU�D�9��>��m��B��"�q\�`�C����GD�`�*S����y]`�ɱ�V7S�{�
����wS_��� ��?�8}x}�
޸>�#��%,wD�v�q�w=��������'w��gO�����I	��W��3�jZzz�Un*�uj����D�����%'}2��\/�w�T��]|r�����
$�%W0�%�.1��3�$�u��1�[�A�k�����x|�k�]�;Eb����z�q�`���O���|\ʆJ��-|Ka��^#`�.j���X�Ĝ2Dd���KA������>0~T�t��ֹ����Fiߍ�30P��Q��v�`έ!���[��13�������
]����Ё�&E�������zH�/dQ�7e�����J�Iz�.�r�@����b�����<i�d;c҆�s�c�_��"��\kj,�BZ����%bz��ZL�����	��V�[`6j�b:0�=8�����NȆi'K�~#�
u�o��i�$�9�G�V��p�܏�Q!#_:��4���)6�*��:!����V���>3�mq����=ta���g��u.�z�全G<	�Wo��U峇��o��&�y�G?	I\l�U?=�����2��\�]�rY=��E�O����z�߂�h9x�}8R��r�]�?�����ㅦ'����j�iv�*�ݔx��1?���L��b.��E݈i@`X��`��5�ms���ȋ��}�I�j����$�M��w{�x�k-bl,`�Mk��	���>�t�&�1఍�y.��J9;?�#ǌi^?�(%I�	����r�Dp#�إ�G8�Y�#����4$%�i�L	��?�Tm���_��H�)��SE4J�*>
�*վ��W$g ���p��C%�+����;c��j�Ean���>��ډt�{g�����-'�0��@@���c$����ё�kz�U�|�R��d�>K�	��.F6��#�XK�g�|�	a�Pn3�(�!/G���lP�ee�Ϻ;5��x�Nx��neaU��~b��u���?�� i�m�~�}�(�v{�x�$iЕY����b�x�D��B�Q0*N/��PL@l��,���7�&��7N>���q��/ߍ��`;�nOd��}56�{e�k��(�/�X��~��u�|�*t��"�ƭv@$'"�~���e1�����/�| }k�kn���+�u�fH�<�R�o���Gt䜣E*�5GZ�_�2/ޛ�D9��2�6�o�0iU��������O�9���ȣW���VC\���բ��(U�4�\�<�o:�l�� W��V?���N0�l�O:����|���?�%��?���1�:ٍ~���%�?��*�Y/|�k�~Xc�x=�� ;T�/�G_Y�|�82Vj�Mg�ߵ���[���$g[u$�Y"��.��J��7tY��Vq��xE@5� *L-1;�O��T&Z�s��9b��;0I�cw��$J�|%%!xoF��;���͕��m�ϥk4����D�."����� Zw�8�~J��!$p�,�!�����\���#/�f�|��N�r�q�\���b$UE�8����o:!<blGI���M7,eX3<��I3��f���w�W�7c�����?%*Z�^�O�Qs�I����	��)�B)|��v/X�����^m͍ȝ܍�2û~Q��q*��Y�q�����O�&��x����}O-��eyq��-��=�}��U����]���t�	�WGл�r��c:Yǁp �����^hz��봜�pY�酜�mbA������Xo1߱��Z�t�������n�����:)}����&�鱿�o�M�t��MSjc�����<�H�_KM�<�B^�Gj.��l�����;����W߇G���:_�����*A�b�S�e>ʝ8����q�Xh2�	H>�ˢ�h{>���[c�q�,����0��5SPX��=��Xj$j�Xd=55ͥ�o�h{��į���Źu�B�F�W&v۬s�uq��:ĪK���\]����,��A	�J&��p���ϒ�8�D�~���̩|GWSf�:�z��>xtc<������*zי�})�)�+/wuYu��h��!�Ꮨ0KW�.H��	s=֍K��������pg4�LR�Y�s�;�~,��z�J%����@������I�
]���y�fE��"�^�hV�t&?���4���Q�bj(�(	
�xŗY~��3�s-�vC�׿km�h�W�s�Q�d�Ӑ��#mf����oU����'¹��V��S����	���1�K�+���O�6u�UWĨ�X�6�݋��ڠ�Ca�l����U,��Ge�G� ��A�ht�X+�[��l�F�V+�HÜ��Xׇ��S%�����������f�׾�x�+L�����s��iV�����{�֨tu�?�aU�!�z��*g�]�vvܢV'�?.v^��n��x�Ē������{9C�ֶ7�H]��Y�h�蓥�1�K��J6{���^Ks���Kt�ڋ�>��?4Td'R�/-��Uk�L2ZIBJ�M0 r��������Q�����3<)�/@�%�D�'K���p�\[;f.Ͼ��*�`;�Å��2G#$���[���	Ys<��"5;Z�Y��lh �ҥ���ѻ����nJ���ZK�����\��᠍(��	��FJ��������a�7M~y�6)�S���Έ@á�h���5t���qB6�6��hF�����\{�4�H7y�P�����>nq���h.1�'��1u%Hz&�P����Ņ+�3+׿����k�I����J�eܐ`�� z�k�F�	�����:���1��8|�-x|�y�Ĥ`\�����h־�g��{Ө�}�7��n�4��w���~�ez�a$�Ӳь[HOX��f��b4��g���ٷk�e��~��u<ϵ�' ���v�B	L������ ����j��,,,4"��sNb$��q��*���{S�wl��[d��&K��o��n�Ȟ�G E��h��䉝V�$^S|:*(��l�6H������i�N�6�[Q+�����;H6���]'�G�N&���=��"l�8&U|��z���S���٣P��q�TJU.|���Ǽ,ỽw�mCTY��[�ӿUB��pd�s�U-���x� o�<���T��?�B�b�5}�_҅�n3�\~NBޝb�0�ի�,#��k[��:{�͒~K�L�Q�Q�$�Z:��~�]{$H�����ǩQ���-լ����cgP��X�HHT�ݪA�讏|E�W�;b���l��E��"}>X؏~�*��l����Iʈ�I6m�r�����g�'�߯Mp�{���@��;�����l�|�K��I����7j�K�$�!�h�cP�.��bE�w���HAx�b'�H��A�eG�,��l�G��z�ӽ�iR�//��؎�~i^����1K*�	�xh�z�A�WJ2ph�C����q��yԖ�~e�F����0ҮxE��)��~x��*:Y��6\�����(��x��q���I��&�X���N��zym�
v�5�苛�zme����*::���f���������e�hn_9B��D�ڞ��n?�8|�{���Δ'1�:�wӏO6E��q	�����Y��~���/ꪯG�����`z��`\�'��
��<�1����^�XN]t��y�գ� �~�'~�\����"�U�qpp��cf���~A�|,(.��YX M����6$����T�/����}���/��=8�tij�iIV��'N�J,���3��	F��LF�V�$��ٟ�b�͒�U10��L��ȟE؍:�z��.�����ǬNe�I�8��A'���ܣ��)�Y.	cR�Ϩ]����s�u��5f�����EAښ����]iiyh�B�pۭ�R���Ѣ���z�ڕ	3����j'��.H��l/d��1^���o�t��p0�2����~�l����(�^d����U����<eY$�Q_��G�: �
'6��,�ٴ���rT� �!����Ά�Q6��_EՎ�KY�}�W�)�R��.��Z��E���#*��#O��B�o�u	Wx�>�ܫ�6��t��^����W@���E��{���Z�}��g"L^���C�b�)%�Kv	.���z��x3yM�>��ۣ���j�F3�0�����	����I\�-p�Ut�'nj����ib�K��@T"���h��Ee�m9l.kC�]$��ی 2��9�g4:�Fp~�GK� �Q���R���)�5�&� 1����9�C%.~5���b�l`����I#M3vY>#��nlgq;�j����	�@u	��. L�",ų��U������e���9�M�hp+�G�g��1��q�$(�h�;��%��G����m�|���c��~���[>Ѫ�O��4Ԟc�WIש;}"��N���fE*�|E~���~e�q�.��}Ҹ��ko���^aq�&מМl
�cYT�I�!)��a�q�f��	�п ��
�sg[Ib�g*-|����*haa���~����G��~)J��]pfv�����-�=ȑ�z��N�?siɭ0�`����d�⻸��T�je�����8G�����^2X������+�%�|�EGH!Μ_�Z @]~-�7�%�/~���Z{zvu?��¨w�� 'C��䶒־�f�����%��4���N������W� �+S ˿.\��_�knu�)1�+bfڞ�W989&�7(��g�NK��7����@d�)�[����\��M�҂s���O?%�֦+?-�]�R?��A�)�i[���=��'��kG��d�V�����ʱ����ۆ��K/����T�Xnj��"�d���C��m �|�.n�-��P1[���@���c����;�B`�g����3�DhAzzU!����R����q ��)��:�{/��F�'����F�@��� �0��:�{C��+c��y�l]&������joѲV#U��e��(%Y��`�s?�W�i��U>�{V�mtG��R�U�O� ല��KM���:�k�)s2qN��ZO��Eh�@�����.��D �kk20��p��}3���67#�u��s ���Cq�@%�U��l�Ω�����s�j���+�~�g�#?w0��jKI@#����e�A�&h�נ&)Ό�A�u��"�X��U���
K|���f55�MW��~�h���ǧ£t��A��Y����m����rS�pX�ǒV�&�h��9�
�5�����s�; ��'�r�=���o�����	���+~��ib*|�:''����E�b����{Z����j0�~����7�=�q&06��q�-��t��}���-�W�s���U׏�g%Z�?2(d�b��N�M4�"����1ʢ�-F[������转"yȓiG����B��my .:kZ�F������&OU�G��,�?��s�X���\Ậ� �݋TB����6о������L�1y�C��kdt�x��V��:}"���@ë���P���h�CKaČ����x�l�[�L�<�� ��o:I����%�CwRLt�$q��	���@Հ�nc�*�[���/%�"Ÿȿ���/�Y��髏E;�Q����+k�F��2X&���U8W�J�-�f�-_��BAc�B���k@�@]��X�e9֋;��c�r69¸�)��T���;g>M��'��:1�a��PcD��+b�w<�&[��7-���Z��%.��(D�A9��e@'��'�a�H0�bj���k`u�Jw�S�H��9޴6w���\W��֥���.'�F���E�8�)�;���b%����R��J􎗥|��6��mD^�p��ى>�Kq'����𹼆K�}r���6��l-]����'��)�|��2��R�j�.8W��nZ�Rŝ�l�]�Q����@�H�H���q*��Ҍ�I�{��rvӝ��kI�I�&��Z�	"�q%I3��w��=��:&��,|n��k9�^1���A³2��?�q��R��*G����1~"9��7��-���H���l�QSc�ت��4<>^�'ջ���ׯ��f�Ϭ�ߓ?�6��;O��@9�������$�y7��K?1Ir��b��]�aěk�7	F.v@�����Z#�3����ߞ2;_��ģ]�ۄ���6U\]0{��77��~̓(x:�����Vv�Z���2rX�Ì��4����F�>�G��Z�p<�5$�3srv/�5k��dʱ�c�\���c�]��;��֗����VII)�`�Rg��	q�����a1��ي�u���y��wQ^���뵪��L���7������BqA�o//�r��������9������|���p�{�tW�uE�%�!_�(Ta��<�>	&�OnBMF�^�u#�RP�ŕo:�6ꢘ��w�^r�?��^oLd�9C0Õ]&�w'�l��P�=�a����r�?>�.v��s�ݻOs=G��H�x�����?Z�]�8�-5��e�&��A*:�O�O����/�.{z~Z��5���S%�3�=ay�i
���T?=�L���J&�ˊ��Y��^�=�k���1�t�o�6�Aos%�%d�˒���?�ӞI%���E���Û7聰�%?t�e�0��g)�	Y�u�+[�R���ƣ�d#á����V\lX��D�=���<9Y��O���'[��m�'*k�KZι�^0�]ӆ\ĉ��4�Xi�&���s�B}���Uj	�V��j�6Y'�wJ4~�:��bq=�wE��C��/Չ�Ҽ��6h��lo)��7;�:���h<kM���~p����Pq���a��T謧Z�/OMW�I4��&�`������O�
�3{��|���װ�:V�������81U�>5Z�؂�-��f�������WBj%���ǩ�C�X&=�c�cqc�褗!���w��}������8k���o����.J�T&��`j�|o�O|��EC��m�C��<�S�)��A�<�`&�D�L�������|$^�����O7�Ã⣺�d	��mv���"��l�V+1��Q��4ӽ���Z[��z�a��/�m��[�LrT�9��R�`�=�	�~�IEy��<j����XQY�_Wg�d�����Cg!�������.�kFLR���$���&q0�c��̾���v{�u6%B�Gz"���'�w�Jv'0�Y1����k�9`i~@�����0H:Q������1f�KC\App�AB[?�T/\i���FP�/���UZn%����uo)���^�=���o��U�?g���� ڞv^���3��� t7c2Az����bR�O�j���͑��js��Bu�򨨳����hO�~cXR��\x����[�����ބQ}�p���OC��Y݊��/�bwQ���r��"dz��c^Q���u��+�*99��n��ߛt�)& l�<��k�W�D�:B�z��Y�vu��x�%2�{C���=�+;[�q���`�^\V��`���m�����R�h�sq(�4D�1��獍�/<jn�ma��ѩm�}~��?���Aϒ�iou���ʊ�߆n��Zhr�R�F5��t;��-.2��m��>Zq<<C�������0L�F��:ZZ_K�o��"�&�@�M釥��W���<�^ڴ�.޺#"�&�ĥ�j	ؐ[����~�"�_��H���a������aG����n��-��Ĕ�^^�e"�a��/��~�YzeC��L��7��Ό^�M
�Ο��$���ϔ�*P������A�̳/"k��ʳ��pp�<�D/�i��H��;c��������O�H��@eq��ϫ�)u��@��lV��w�����0�z���U�EX��7�`p�~Y�L���r/�z���\m+W�*��W�H���� ���	``Ik�LlmL㕢5�/��D�R,���s
:H��0�?�}��O�dw�KA�X4*at�*@���5�>(���Y�S�"yx��Nl�c˞�ZA��z��W�Z���U���h��όٽװ�^��-`��>���B�Ha��wtT%Q�g�6j�N���� �w�r�}��GE���K��
t���=�2�$o�xĈkX��8<�X��[���^�u:Z�{P] u:7mˇ�{4���"�B��������i�ҝ�Ajlвl'��+����߻�x�7���8��e}1G�����bO�)��k�(�}�;t
���`�3{f�go����BJ���ƤP'�J򔽴���5+&^?�s����Mnp@ܟN��U�������Gm�J�O���ۡ�7~,�`��h�ݹc��!����Y682��쥽�2��6�F'<y�X��"�%��[~(���h&�;x���H���.������L��U��b�3~���e�rj�S���s�@6����i��V߳�#���!��"Y��h?a*��?�hz���W����{�el�������;2Z� � ��;�[�
oT/�9�	�j6�ڬ�/Tڈ$��"@��?���7�)�6�K�@:������L�i-�;���>�q5���Gl �����rq9A(J�;z��*ˬ��f|��vT���m��'��X�16��§>�"�}Tٗ�[>�eԉ�=�Y�_zK��e��3p���;���k`G�L�y�@f�O���U����AA�~���ی��-�3ӡوS�/���v�VE����`��	�
%e�'���xى�UKg����>V>4�%؂��,yH9/�]n��(('�}P���{��̶�d3
��c�TfM��8�AA��*Х^V��E�¹䒄
�(ol#�g��CԵ�M���������l�כ����bԺ?;��X�V��/kO��t։ ��'�xcy#���s��3�-19��(�Yt���c� ��W')�&��	�Q�B��jC�V���ۣA��sA%�&�P%�t�6��Â'��:D��ĉ��M˽q����->��P�#:���1�e�[�C�94��_f%��WU���;�֗0_�Dkc�_��|2�����u�9psWx����;�Blj�r�fe*�~� �x��>�J��Ŋ�=��	�ˬd\���)�֬�*�Q!x"K��_Jְ�F��~�$��J-�}�U�:_gc ~H�`�` E��:����P�0#w�͞�M���0��V�|2�ҏ���РL�З7�w��>�1qq�bno^@��x�ѥ�9S��UB[m�Z<����	��Z�(O����Z �0]˝� 3wc�6uZ�]�&�J��x觽��l�V�u��F`�[T	�/��H.e�Mu��[#�Ӱ��|��}9�:�O��^����2KUW,��Zn�\=����,d*���V�0�4FH���h)�Q�ńE־�ș)��z�����8B�a���g��~��
�E����jD}d�L3z �P��ed3q�"V@ ��M�I�P|\�bH�dۢ�&sp���
�_��(>����+�A!]fa�Y$ߛ
���]o�����C�!Qy{,�T�#��v�S
��0m�KL��c���L�ٱ&�+)��>JʂL�w��
���:�N��{��_��+�{%.���5K�8���gPn��6�SMz��xM�bO��l���ή򍙈t�>�hb[��Z�N����6�L��֘Hvo����#���A�۵�K�'[�)��_k-�����y_+���UX��0x�pYGk.��j4�X(��3ګ�0�)2�t��d�
�>n?�x^}'��I��qe�m�o�df��U���V@�Z�ʼ�(�*�]�)Z��L���]Y�X��0��J���劉�����ixy��������@8����R�ʮ��]�x��Q;t��p��F3����jnU����E
�~��kL_�gxW�{yB����'��WW�L���H��¥[e���\�c7_l���L|놌_���`S�p%2`�+�QLR�R*����a������7U�M|C�Z�+	L��le�CJ��5tL��t�Ҟ�#�g��3;?yq�t�s$	7�u������&�.���s]F����%���*�tn�X�j���<�^����|�{�7��VHm�E*��|T	�����>�1�����r�o9�d�h��5wl��o}XQ��F��MS�ה@/G�ϊ�(*D!����w4��X m��CA�Tk��|�N�`���\����VѸ�~^��f���w�� ��w��H�,��w���h�=H���N@fAg
���hp�-̕"y�+��8Dr�.]�(t�Z-����[a'�����2Rod�̡UŌ��d�hVCs?���~�gV�w�G��n}�@J*�K�M�;�H�e8C�	��\T[�����uI?i��G�u�C���C2J��R��ǡdg�]F�ٛC�E��=r�^YgSdd;��l粝q�������<<>��~�_��z����޲�.w�ͱ.?�ߦ�׶�3T����J6J0�*M�9�}+��{�����/�W&;�5)�Ѓ�3�'�#���:��j��մ~�V��e� �zh����z	4�_yO�\)Vk��r:|ڮy)�m�g��;8i�R"Ч�� �o����E,�_���\�6}��\^V���bnBq�����ڱ���u%��X5�~��8B.�+f�q]1�D/���p1ۣ/7��p/�}nñ���J�v�X��3��:\�=b�L�?�Gl<W��v�Yk��n�O�^��.p��A D�U��?��<�l�j]톷hn�۩��A����Wl��׭7Q����0-�v�v�+�%p��Gc�i����?�v���� �J��1� &�#G 2�T#�Hܦ٫#���E��6݋��' ��Wa�����;�����u@��҃+��Ư�|�9Kǉ�>i��)�,�5�V�\�����`��b��}�7򮑻���
m�\�{2>Y�	Ǧ�e��?���y+#u��⳥��?&�*��ԪS�w<�����)DBL�.)�$��_�M�)�jШ\��y?����}A_�dD�^�	}AU�i9���]L��>Ф��3����?�	���RT�����r���$ɭ�1�t*ʩض�F@~��m[`��ע���i��c��?sn%L*x�}q��X��I��ծqd��I����cg�<�`�B����̪q	4�	�5��(����9������7�>���]���Y�c?S�U�u?BI�VU�N�_Y綎ĭV�z�6�cZ�HӤ���>���?K��D�`���D�n~�y��Ѥ��DR��%�5(\0!��ɘƥ\ȋY�e9&�&`Yo'DD�+��`Pg-):��TNi:i����Ҹ��ީ�1�);z�EF(��q�c�S2'����v�~���n*�^���<��a^Q�q�>��ܫ�K��F}<�1��{���s���!یWG�[c�Q�
�	�\zTKk���9;`�ACZ�Fq-<�ҕz�R�z�y�ag/}yd&����-�f)'�U�6w��3ß-��Ǔu�C���oz���'$�F�P�΍�aݲPk_O���@�� r?8Ֆ� �Eh�42��N�w��
��4���{��1�&i9�O[���0+ݺ92�x�p��E3��2/���eL	�� '�3��lzXC�{޼����b+R��^Z������2 6^2�
�˹���^]xp����i.Ñ�f�&(���Fc{��2�꘽��hÌ��G��@QM�*����B�<�a�q��R�`��nN�,
��������c�A�êS�e�e�+�@��S���f�c���H�nr�+T�<!Q���2��{��e��$4��F�3��Jy��G޲�h�7_��u���b�}X�
1��mE2�\?����`&���?ZN�H=�|;�3/��q�����rS}q��GW[T�?����� ��I�6�B�ō�!/VW�;#T����3���,z�b ���)���8�ڗ���sw���F��Sj�%�o��//�0 F���Y*g�H=,$u��E��g��������j�Xwu���rAS�f7R'i�3>@d��k[όҸ��������r���e�|��7~ߕ�����[��:0�x7w��ϊ��b��;�y砶���!K��i�bY���n�7�.F���"�#o"���ʆ�Ў��C�ޱ��SRi+ƸC��kW x84_I���ǘ����a����������%�4�jO�5��~��<5gC>:ec�zUI�&-G�и 5�sJU�<eɕ����j�;<�����g�[#ys8���������gu����0����꺣��ҷP���4^2�<�Dg�����y$��dCbRm0��h�������S����:�5q�ϒ��b%���C��w}%�7�v��_��	���g��y�k�/��RA�����"���)�0� ����d�b0E劷J��;�Pt�����#:�΂����)(p
���
���\P2�+_+�b�4��-���Uv]uUE��5a �]��a�n�ǋLi\q�d����ڵ�B�)5��_�Z���[�ҝ��lP�J���+�]XYxz����������c�e��ɪ��9L�ZM�l�q�!���wz�	�<��I�VT�h��9<^Rx:l�(������\鮁\J
{��r�z��\�n1�*�� ���_�"H�i0�*[I�3��Z�I-�Ix�Ys*���%��D@�:!j:��k�͵B"��(a��Ѥ��[��=`/�E��m�� ,�2���H�s�N/X�S�ܦ�x�2�kM�m�'�_^e.�q��uX$�s����������S���Fb� ���wu�M7�7>�Tv�?���i���Y��sp���s�K��O���q(F(i}�m,&���Yp��4v�s�
�7=EA���--��ZL���O$Pbw���I��S�:��~���Z��{�Y�6lT7����lF>a��7�~R��Ư�4KK�WV����5��Evd��U%����Em/����P�M�뾆� ��\��~�>ҕ������ܞ�87!�:-� uHqC�R�sד��ƺ�}��j�7�B\�{^p�êwgX;\�y/u�)�Ťu7[8�΂�@��/�~j%��j�t,���k8	p��Vwww/�)���V�����C[����tQ�:�����Qlh��̍���rr�:;&}���+�Z���N�v֝��O��KI��D�����}%��@|R��y�|���6�66+��6i^c���� (�Q�Jle�]���m948�g�	Z�YT�(�ԃ�+�w*�٣��+���n�&D9͋y����Lfj%��*����%��0ҌXިs��Թ���J���8�p�ɱ�徉�jpS����1���Hzaw7�CF[��uΈ�e��0��]�ė�2߿G��5�L.�1�48n	�c1YB�02	�V�.���0���z*`y�a�?[Ɨ���דB���t���AN�{������ �	,u�|@�Ic��v�v[���&f�=t� "s@����g�R�rω�"S2>��*��`_�g�Ғ6N��d�2ӛ�ܵ�ɾ������'����6�ɖ�OV7<� U�׻�d�OM#xI؞%�e�ɂ�
�����m]'cW���������oFRcۇ�������q ��Ր4:��<V�]��Mq����D\ĸq�oM ��פ 7�t"���]vzr�Y�ٍbsJ56����~u����v���t��ٲ�݊J�n��������T2��![+]]����.i��ӰQw`/ԍ��y�+����+\�J�s���u����#���M_����@G6�륮��b�'�0؆R���+��/ǩ��`���i���^�8��'b\ξ��^a���3�U� ��W��T�O��.y�����Jq�Kɂ�k�����f�j/��ܵsr�U4��p����g�
�G�U:A��ܒP���+4grj�t	$�U�D�Z~���;O��c�\\ɪ�tnj����Ozv�§���h3!=�a�~�-��X�g�p+���x�f��p��G蹕��=^���Cz�.�����G��§l`E�^���e)�����D�zD͔���2n��dkòx��hfG�?��/�9��1�cS_�>��PǹzN��5�ׁ��Tޢ�E�X���'�(Ү�PG� �T !��q������	�g=�j���&��1�Y�2��d7��L4��� 	?/�J�{��Q;P\&��/������&b�J�-�q���f�zz3�v|�OQT~d��Sy�����hg �X��cM�pt�4�a��� ��?$MI��T:���x��OV��5�Q�/��?F���q�8��������}v�4����A�:�䍱��ÞtFo~8c5#9�E�%�D�?E���wU.�0�$�6��MP���݋�iN��hJ|�CV������h����U�s�^��H��F�ݷZ��|��w�Y ]
�������Q�e-f�B�Qq5Wk��JkKG�~TY��wR�{<����TX�h�Q9�N�����0"%�5�ʪ�My������8=]r�5�S�|��]��Jf^��;2	�?�j���y��к;�x�"������-B��f��0e���lgNNL�*-{tܛ6�_�:��b��&ӱ)�t�1!�`�5+�Ǔ��%2R��K�v�������>u�K!Ca����K�b�WI��w�����ib����o���4�lS�qq���U�Ya��Wɹ�E��:���k�Mպ���'#cK��Ι�SS�f$�h��Y�G����Pc�ڞ$wT����`�9�W��K�%͔<�Mã2{%����!�3�FΟ��ח�̒�-+ns	��Ş���@�����I{"6YC�ΩU�A�O�jrf�rrzdOw��b�9q����#OJ 3,F�59ri���М���?�����'��`C=�9�<��� ���3� �_C�e�k�_#3�G>+)��ת�_LI\@�
E��kKx��Zyڹ��&���D�J�,ڑ���H1��	G��C?	��
ZZL�M�5�:���A�H��r�y
�ic5��FX�v���f�����*a���X�=�@9��s��u���q[�2��9��b���a���Z��5A���&���+\UT{t��Ԑ��T�ܕ�����q���,���ʎ<���c��#�ڤs���F�mw�O���/��G"Q�w�Kv\�
^o_~�۷^J[�+�ze6�u	�
R�?�F8��h��U �5-�lT�jvv��}C�ق�Wh�f�Ŗ;h8���D����L����ޒ뉂��,.6�`�I����x�/}g<�(a��q[?Y'��O����
�*Lw�e�ySL��6���{�kwE��2&�v/�7Xʁ�RU/1�;�-�e����\`����fve��B& 3<��c�N��f���g��������k��`�GM�N$k�?n�_�
�X0?��d�� ;=�ϧ,q�y�:��*�K_�y�QV6A"m*"�������N<\EWhF��!(u�Rv�#�T{dE	�Q�1'��|�>�z� 越:؛w�#�[2�����B'VK=�<�	�u�
����ܯ�|�k�v�ڄ��u;�b"�җ�����@w��f��Q����eee���IM�H�e������P��S��e9�j��g�^��|t�f��]�
>���9�E��w쮫a���W���2���?:-]�R�-��y�E5{ś�ǅ��7<��%Z3Nq����a'�	�*�
�I�UK}�eu���C8W�p���C�ݷ�Gd6k������|6���Y��g�%ZU@;���Ez�29�Hh�d���Ɩ���T��i���������G��kT�k��D"-�\}CV���j�wh*#0#�~nX.b� �m�^*ڊo=�^�kv�&���G?���@
�h�k$h�o�?�\��ɃL���M7�_��c������WI}���C���&&�ʗMM}U�0�L��B2TJ����9ܩ�cN5w�$�\�F V�;8�ᮼa�m�����M�r����G���v蝽3�t� ��+�o?΃��4����"��e8;exaQ��e;7�@Oz��$�wd|��K��.#�twk��;��|��::�~�?C�����;R��<]۫�bu|�3��3=�c��*?�hvwLFĭ
T��Q�а�����������#;褺�uD܉�Fo��٭l\���Ho>j�P�Q��o���類��`����N���v�c�����bg7��Er�M��L�i��7�9�¹Ju?���3����>��G�D�1��U����oG���hg�\B�n�Oԭx��Y���.{�!��̹k��/;�������G��E�m�Hd���E2���������>up�I�)}�8|�ʥON~�n�[�h2_�l�R�VFkP%��G2 01���?�8-�+��0�J�`��ѕu8��T���H���1Fa�o�������2@��M5���j9�5�HW�G��"�vn��~0�sv�עe��K_�[�� ��Yv�5��*̤���8Kdd�p�,=#L�q��BE3	ܳ����t�;/юM�Y�Q�O8�yy���.R�������e�T^[�?4���GUuOɗ�;����;vX��
訴hl��1l�7��ß��)V�C��R�i�7�v���&7z����s���2��y��xB�E���;����^KYډ�W<W��䮘ߕ0����M��`~����x=Q�$U��s�;⨖3zuW1SF� ����NMSC"ā�� 1�C�K ����O!Q ���A�H��6t<���o��4����+x.���O��>�����w��i�� £�m��JѾ����7�T�^%oiکH� �j�l�JIn����q.(�ԍ�[#������q@���ud�]�p���w*ë7����;�;�b�#S(�2��{p���{-Xv�f�[�-���a[��.�ҥ�ub{xH!���(hå�Emu�'���-���5�|@�9/M�0H�Z���L��wzT;=j?.b�0$+Ǖ��jњOkw�
}����!�H�n��(���n��5�>#q����m̯�5H���i�V(���=;�u|�4�n߹	ݤl�e���,b�cW�laZ�F ���R�2� SO��s��3_����@ ay�i�x"��xzz�ߨ�
O�-H^c���c�>�B�����J�G�w(\Kߖ���*�{�t3�:���Br%�dx8a`���mq3�x+ڜ�A�봮�xf�X,)��+���L��[UU��M�����y��{�,^����Jr��}rjO<�z�>!;z�L[[�.�~n_	��٢�ܴ�m�s�#p�*lu������ũ,^T|HV=f�֌|��cR��Ep_q�q1\�_�U���)E'���9����������Q���b-��ט���]����t_�����]2h��7���99��V��C��b����	�F'��:�|���[s��v}���w��
�x(P���%t�O�(e =zW�1݌j�2�d�.(�_,�6���56�۷�K�rk�$o��vK���_bR	�oT�W1�����U���Ȭ�BZ�u�P�avSp�
�9F�:��:��x�K�d �"a�"}LEҽ���pV㙊x)6S�k�p��K�JJ��1�U������#㛔,0>k����h��@0U�]��L=���k���D#6E�ȸ��;�59u���|�)^�!6�U?��B�E�i������=b�]��L����L��|�Z�[�����_zg(@���{=Z��a;O�*�`��q.y`����J2��9�L%8�*j����$C�b�o�ܢ>'��74���6A���u�*s�"��bv���C�j���K�If��R׷	�8r�����j�G�+�����"�?	���v_�2��*N��"�<�u��G���ok��R'��&�����N��������Z��ۢ"mm��'�����r��*����Ӌ�eN@_8�
����8�p7���Q�E����z<u�m��c|������*��\B�v������b��IZ���LFT�Pb}����z���?�� ���Zf��x\���_A���@���Z��%k݊2�ob(^,�`hO�58nK
>�c�@��ż��`կ��!���rU$K7�R��z��O��5rm��OE�Q���y�s��ϛi%URf%����ƕ��?�o��B�c턻��Z�O��K��g�gt�/�� x �\5�^�JK�?߯��%8c�D������yTK�����k�Jis�/�Ѧ|�T��Fx?�C$�����?�������T�Qg�(��u�������o��%O�c��	�(�;$�������)�v/�,	��/s��lṦ�v���Jaa��[)5c�ԉzˢ�2S�1�N/��6х���A;��X��o�(k�1�~�8��K������ԭa�?�g|րF���_�������+�!g���99=�	lt�
:4� GGzG���[��῁��I���^z:GQ5 qLzT_��4����q�V�>����M4�ƽ^S�̮�A�p�a��4Dj7n���{���_F����x��PQ}s�ݻx� u�_3�nk�*�m�g|�Zh�xA����M׍t�?9��O��.�͕�r�ZC��N[f���t���sХM�!YJOV�ܖ��*"#:l�����i�*�y@,.���1LQ�92���86� �3O�YQ�8Ε�%���R�#����/"�#Y/�4<���%W��w�짏_��:9:t� tI�-(
8|ۺ���{��b�P�i�;]�:�6�)w.�W:�K =�'�E:Ml���T��P��4�1Ǵ;���z���^~�
E��zܳT�������X�T��t))��Ñ����:�}?�[�U�:�K����qg�pB����~L��bBl1/9@
`�=
���C�:zc](ֹ���q�CQ�hK}�C"��wO?��'/��1U���>>p-����d���iSܾ	�=Ɍ�#L�{�bzZd�U����y��ŕO�'�P����c"NX����P3�[�0����a1՘�/�$���
��2O))i~V��Mo��6-���0�����F�-K?��<=k .��:�t�8s�U�h�?,5�n8��B��aU�%�Mv�뫗�ZZ��Su�6h�+L����/����u�2I������u����t"�wx���Eh��*�u������jn�G���Ŷ����/}@c2���N|��1t��������Q��٪!�wi�y��^:B�΢�r�A���}h]740*��*����o!������u@�Q��D��s�aKc3T�a�|�9��偁�����E�6�ǀ���vW�Us�Ne!mb���g���z��(�|���]qU�I��+������dC- � ����D4"����F����L`z��1������umA���XX���{���p��,r�n�~�9Q�^��W˲��cn?��z��O��nfH7��6��� |M�maQ娎��I�n�&��hfL4I��>�r��q���f��_��A�/. V-��D�zM��᱇~|N�ખ��^~�a�f�#7�B<�i��y)��򦈕�&D�C�ZZ)�j[ ��"�/�U��|�������ݲ���gE���9xj��O�b6w�s��')����9������E��d��|鄔���%���s�'Vk	>;�z�)�0�8i��O^��Mk���I ��T+k�
uw���0�6X��Cp����މY=<٪����cJ �f��xU��~�F))W��>�ы��s�v���V��pK�����m�A�rrچ{;�Q$Rv3���콖J�O�Ύ)h�0V�V$�vl"����L\�,��nUSK���h?��Y���pI	$,G�38��o[�������j���*�7*�L�_��:�@6��6[hՔ:��4V ^a���!U�[j2��Qǭ����=#����d'S[>2D%��-Q֧��'~;��0"z�W�DbTŊe�5��	R�l�DNn�v@!���)��,7+���*pȅ��]��S�����E��Џ��@��;��)J��(�aRP�����b=�ֻ톬�\ն.&PӀ��d��_/&�ج���q�!�pT�������P�`F��C������c@�
�N�7�z������V/=K��N�I�u����͹��h�������r��N�|f'�3�e�>L6km�O4߻5 V�u���Ϥ�w�Gud����Oj+�������ߕ�*$(��!��ٮ5	�C�z� �U��v�5? ^���yd:!�x<��c�@_���Y���97�J$�����On8�0|� `��L?�-(��rÁՍ"ΞpR�<
�B����V?�}�ъ��A����\A)\V;���aDl�%p�,�e��\ D4���H��!rff�����p��^Ydʄ��F�<��w�ܹ����s&�R9U��E�Y11�| Fr@V��R�#Sy+�^��J�6�V`�&�S=��D� S�-��;5�w$�Zd�;Cv�i�9��2�Dԁ�ZFI=.Z\�{�^�g4y��KZFZ����:�6��e��j��Q��W<��w��B;�J�8�������Wu}��,R|��K��?3?�xc;��ZWn?����\6f�JM�N��f����G����d��!Ƹ�|�5A羼7��᪂�V��L�\)u��^�E�:�vڤZ���=_���PN�h�o�_�)�o�Ç��/�T�㶑u׈��ۄ��o n;t�T9�����{�^�I�(USUU�����y�}?��6��m�nGJ�~����oN��'�U���v �5N��uk��Y|��i_����b=0�y�D�{쎌#s�K�kA<.aжv�g�N� ����UBs�5�5O�� ,��>�,�Oؓ�=���#(����FM�c��H�A�=zm�m��w�Dj~^��ܢ%�6g�|:�SW�)���Ç�?�3�\� �IY0_��goyʙ$:�C� �(��ŗ�,e!���۲@#6RX��?��/S��|�`�;�Ƅ#[��5�����k��f�P�Y��s!L�I|V��UZ������E:�!9FuW�]=��^:$��?�h_�ܼ��i�=|fF�^�J6�jNlkgp],�8�yL�����I{�`�j�%ބ�q0�٨;� "���.NFQ�� �~�"tc����Cᛲ�1S_��R�ƝS�����,�R+|��y�?�;�\����ۭg(����\jn��C�X��"��Q����K���`�K�-�÷6��������."�}h����υ�5� 9�`"�9���/�D���xܒ����+3��"�Z~�o:p;�~�(�ҕ^@�QS�*A��:*h`E�\������(��.X�L��_;����Т���ܩ���P��$��_khY4K���k��6	9S�e��R���?O�8�,�����H���L�+_��A���a�,}4������$c��ݬ<��·u�pdn�8t`��}2a}Z���zPv
��H0����֘����x����>I��R8j
~�_X�|��R���FdQE72o�0pģ�+�"�<�0t&IW״9��-�tC:���T޶�5A�Sؙb\񔣿-�S41��Nmek_��OmY��Y�x+��A̒I��*ؚ��뜞5�p2�?��T�-�����τ����,=�|��4ME'�^�{���X��VS�E]��7C_d���1H?&	��)W+�|�|lh���N�s�?�9n?3���+���Ã�J.�&"���ǀ$��ȱ��c�/�Cߞ�y�VRm�آ�f�ܟ6x��z�
J5������PËo������@��)u7#��}C�r��9w�?���S��ݽ�8��q�����yT�XLH������5������#>A���/|f����8�6{{N����o�DM8�����H/k�rL���8��Z)+C�����Ѧ&�j��/tj����S߿�Z���M�A���YSF׽��
��#i�ٜ�T�)�wG�4��+�?|=�?�{Ɵ��4C�i��o/�4��-4��0V7�:(��B� �lQ�kR���}��my�t� �E���UW��x�C��\Z�h����ߊl+<;�b��ů�M�%�?Zm�h�]^�q��YM�/��������a-��G�ώ*�@'�]Gto{#�AQWσ-�����ίͷ.9���� (Ψ�pr�����J�ާ�c���!�cl���??)���Q�=��-�Z:3�l�Z�1F7�O�`�T�_L��m��%�.�Qoiu% ����k�_N����ݑѰq�.���,��;a0.�w>/��@�C#w���^R��ԣ�OCq�b�����xg��%� +�@�:#��<�[�(ePyq���Qjֿ�;-M�:N�"P�������ќ�+��T���y��+R��3��:u/iQޟ"g�z�����w;|)K$x�Il����9C��O�-�HK=ه�Z���;V�""���j��������k{���#�%���2%:�{� )lex}�Z��Vq��c@�$�.�/�h�mhP94
=� $yՙY�h"_��s���[�V���<�z�+c� ��֩(w���}�����]�ٙuLG�Ni���~]���(�E�m~0�[�B�p�0E��!�FS�_��>�V 7!~�5b�����{O�A�bgg��+s�Ƞ�NI���
��n9\9AO�I4��TX�7~(^k
3�r����.�F�y��lӇb.��H�mE�U�z��~ooR���o��e����3e+�ދ�I��G�oT����\}^<��, ��~�A����@Q6'2��2���O��W�9$_�wά��/4"���`��8��l���(�b�m�ɪ���d7�)Ӫy�"(�x�"7�.�~�v��ݽ���:�I1H���ۆ*dM�����Pj>���F�vك9r*�����=+�����2���g��n�����JA*aruρ�GJ "lV$�YXD�ۻ�]\�$k/}�ﯥ��w���ɭӹ���(5�(>:8W#4��4�b�J��p�ݒ2�++�*WaVE��6=b�+�yc
}�r8�ub�f��n~廹�zNf�i�j$��Р���AU��&��IC��͂�{j��iM��u@���v+��Z�D�<�k,KoX>�+� � �h�1�hv��/��9�<�H#���`���y�('�Zn��S�?3�gi���gdtǐ������D%%�T5�*'�[�0��$����~�j�>E�ü�nF'�������س�wf���}�IM�]0���O���@U;�@�K��q�D�\���{����k��������ٝ@!��ڼ�F��_���U"SB�4[19��������l�����Ѹ�r(O����NN��}���ylv���ܲw�C�(�}ۛ0L26"J��q�F r���o�K��.5��=N��g-s������qh�߈���.�w҆����EUugמN�>ޟ��඘�vPP�����$��Ar^.�|ە��cX�FM"���'hUw����߇�e�`_�o��O[m�Ry�md_d>'���{I��I��ĺqVɱVQ������7]7�/�x}��ﭪ�!���ʙ6����ؠ����u���)�Y۴�i��$�?��	I��5� R��}dj'���Ĉ���Xo��_��z�b�[��j�ģ���D[GH�`���.�d��C�,�F7�mc�s��,p�L�-#\|�H�TO�7�sT�	��+�3��򩣲w4�� �6�	���"��~�h������C�ҙ�_-JeeK��6�>�@���2IU���2����{��G��m���k"��F�O[�"Rll���+nY�%�UB��fW�<̱zA�p���	���ߧ&��h�J�U���x�>5����mX�Q�Ao��W^�bZ#�fݳ�JZ/��m*ӏQ�%�l|
�B:�����]���s���OMM�ަ���^�gP���׬{��,�dE�~�,|�)}r��<��E[WՆT�^�t��o�A5�yp�`�)vf�^���r\�%n��8����[�k�-"���R���w#�6��9��*��n�I����N{::��v��RW"��ޥ~i]Jr�6fZ��c��ɧ*�����1�?\�$JaR�s�d�8*]�!�ԣ�
���.� �
QHH��u.=��r[Ve��X�<��V��������N;�C�Pk`Q݊J���J��Vrٌ|�'8x�>��5�mE��L�t����c�&�v���R�'R�� '�IN'/��Lh���r壗��b�8H�+�*e3v�(� ;�����*$�[a�\�@��:����Ӏ���J��?��R3w���`��TV����hƿ��9��>jY�Keh6�۰Aʪ6���i�&��[ϼ�G�l�'N%v_)��^H6��s'�ҟ�#!��֯�}�vR!d>���ދQ�ɧ�p���句����a+�?������?���5��ܼh'܍��������XT*�{�����&��R�$STaЀWFTA�af	P��"�N؛G��/߭?�� �t,~���im\g�ϟΒ؞̖�����R	���/�sE�j�q�]�9�Z/3I����
��~QMjj�c�����e���7Aj��N@ $�aXELYU�Ȣa=�d�	���/�c
p����i"�Ӯ^3g���fUCv(i��zf!��!x�y����hwhqG������xNi����8��
>��n��Ğ�*.�9ۡ��uS͘��+OPح��1T�5������wԞ�^~����w����l�O�����o�<Ғz�Z��n�ֳ)��ΌlW��D?c�-�������X30՝NDDJ�!W��9���Q��L���F&:�����ζn��A$�'�r��6e�~W�2���fߴ��� ��;JUT�1���t�,l �jqp�&.��3��qM9{�c0�9nȇ�F��G!�X���;�+"|����z%�(�I�P������O���i�ݞ_Q�H����t��2D4E_��v0l<���~���.���F1����4(�;�.�am�{�IY�2LR��]����ܕ�	@j? �C� �k����4���,5O�,�%�I�O�h�`9�`�tS�n��ouﾅLVp���姽�1/Q_�����*����َ�_��;/��k�u�]��= ��L�y
���m��v@���*�RTN�����jB����@�ԋ�W�դͳhiS�,l�����
�+��C,��0Z������J,�����e@�����|y2������u�U5D�(M��z=#���ck�ìp&�na�ɵ���@�n��f�eA�%ڻc�����n�Mj^��둘+�˒���F���R�~��-��N���X3��/C��MS�e�k)��J���4#��gB?v&Od���2�h�޵e3;8�=�po��Ta������/.��q����N����ߚ�X��7>��Lŏ���p}[�ǉs~�d��g9�¨�@Қ���:��ج��`��d-�W����oV�=��B俞{�5#hPmV��a��~��y���G�rb�������s��&p8|�,�c�"�Lϫ�8z#�Iɋ�ΐu8`1�[�tb$����r��~�
t�|ax��*�V���_�Y53K}���~%(��~`�w����.��_P[J���d��VĂug�qa1Mqw���."�r�7Q�2n�����p.�n=M͎��߱tư�+IU��qg����n��>�Vgb=j�֡v �?�i���YG+�]8��;�LδW�ח�>t�]bD���(h �]b :C)�1�4P_��r/'���tܞ�	�Zρf�d>^D5���q���Z����_����P�T�m��i���vn�=`��Q�c��v�pGc�"���*ۈ�9H������jS2��q�(���4�A�'+P[������F�S%Pͅ���.`�i8I@ʙ{��EVk;?C���J�lZ��X��<��d97sRO Uv��<t��O��	���BvW�w߾���8C�Na����H|�}��/5��>��f�4�ϫi�)��cWbM�cf!-��C]s��w'�yN��#�mJ%S�� :`�L�߈���f5�h`S>��Z6P���-���|�qT�{� ��ҏ�-�2�z�z�M�sf�O@{n��r���C�o=A�-��Q��`���l��\�>�s\�s�9/�%��8äG:o?��mC���[#�?�yp�&(H֊��mz�Dsj�[�#��MOj`#:�m^�l��K������Rd�0:U9�x��H�q%2��.' %=�g�̱��7'Z��uH���Oν�֦�N<<*~<��:9�`���S��n�\Z��1�s4
�슫� ��>�)���o����9����n���34��M�u�#��^#fc��H��6� ����L]�{����(���M���ΰdy4I?��v��Ee}��m��7g�w�c�ˋ�_�����V��b���>:6 ��T��Sf�93�,:#(��\���mdd+ȹZ���:�)O��ڙ�M��&4;�H����5���*L�A��#m��N��� �1��B��q�;��t'��J�w�����͵M�ϟ�$��[�z3)���Um�hzd�5��0� 2���If��7~x"�Dx�Fa}T��V��f�<��"qo��tVpK�p�fP�ao�x�!j�S��`�0���)͵�ī
w�兆7��tT�{l��-����Yr�և_3�'f��p\�W��:�-��b��C"�lP�3�CD�x� ZЧ�˽��⪫��m;v������fa�&W	Q�	���?�����7��<�Cb�	G}�%�v�@�t;�F�W��6���]_5µ�K!) P�8���YM.F�7�e�M�p賿���4᭞İH�N!�b��]qc�	�����J����5Z��AV�����&&iV�C�k�,F:"�i�)Cѳ�	��B�:(�]�T���6�]�}mz�����������~�����������e��l�p��&Wɦ���3�W�?�4�M���h���^�)�?Cs�^�%o��45����\B!�S4�s��&B��EfF͹s�#�Em�����R�ޟnx�gi��RAm�3xƨE:4�-|��־���mIV��Ѱ��tײ���ӥ����N����,g���Sb���cO>��.�۬C��KyГY7m:����jzyގr��
*E@D�.H/��t��Ez	E:!��� U���;�=(H�D:H'������������	[fgg�gvv��99`��)�d��1���u�ίG�9r��	 ��ɩز&e��������خ}���G�w�Tr1�(����%>����x!������.(�E�$r��l]�G>��w�^�0'[�nU��ĖV����E�J�-��P'� ��]g��1�c����L6ED4=���
��~�ݥg"�F� B6ڀss�'ǪX�������&
Joy�?o��Vb��������۠��i��k
�%�&i���k,:��Muƹ�#���=�.�Sں!���������$�fd�8e�1FKǁ��eU~׮
�d���Y7P�� ��1�ך�O��,(���R6��ߔ5/<M���&�I|����|,#z��s�����l�Tqi����Êa�Ac������gϿ��q��F�*���^�%�j�kx�򱠉���~���������^mx��k����d2�b�LC��Vіzoh�*���"GMQA�������B��YI<m !�弫e$�4���w!�� :���#��(m/�>UG�Sl���[:jnpA�]*����.���6_���z
�.���
�w�=ozZ��ы��9u|�Bz�?q�z���4��*��<��)�|fns.����������b�9s���L2�;�l� 5<E𪨬\��d${#A��`��Z^b�����u�lS�OA�F�*�-���z��KWF��w� {�����\ �J!H)�x}9��HE�.�����pT�*�c��3;w��CTd����1؟f()��Z��I�[j���mհ�z.T�o��Q~�&gVr�PQ�� x����F���
͜c�U�����]�Bs�����,A�t	ʶ6�P�;�Z�Ż<+ި[�T��_>�R�\[���2vI7�]�R5M�������8ɉ��r�f|�5����z���&�*9���B����_���3`D����4b��#���Y��dmwK���A�,�Ế:���O��-��d*��Xz�  /K
���?DՔS�W9�;맊Ô�:W���Eeʶ%r�wb:{C:���u��(1y��B�V��^��\�p��J�,[�h&�4y ���h��~�F��w�\�p� {��W���f����]�(a������v�<+ſyϾ)(*!����OKW,�~Wf�z�t^Չ���(��Uk������<ԟ���G�͹��`a�� �5\P��P4��OwS�T���|\��Xx�E.�:�=K�������y�c�1
Y�$c�ο9�Xq�_X�kn���ԣE�/�9؛��%�@-_��^�D+�lG�m�[�d��P��uF��&����
�H�r�DrG]/�f�﨤�`#�$�j����}�<���.�ֽ��p��58���=l11
����T]��,�
���prM~��m����d`y&>��O��^zwM"?�;�z*��"%gmG�ݘٯ�ו�v������RV�TZUY� �������� ���6X�iQ�a��E+�oY$4ߥ�ٽ�����t�wT	s���ʙ~���ZE_�v���¼�Mʨ<����:SY�3K��BSlnM�U��|l��ͺ�Iǀ.c	`�I��r�&f�.�R" [�.y\\���/�K���Vʥ8����I��I�}��=g9W
v��\g�i� J*����ܹC~�W�n��e��}9&���̀�)ǅ(�`/�˳�+�9����n����O�zn���k\h�8\�~9��w�+6����NA�r.dA������Y����o����Hv���-h�4�[ccG��Y|�1]�ZT��T���v?�o��3��mc�f�J�N�)2��r�9�<b@`�|#)1�$��.d�w���  1LKG��I�KA����W������ւ�S�ѫ��h���?���3�{	Ybì�ʞe(�8�o(�L*-H�~��?u|Ė,C�C�t���J��dL#t'CMץ�T;5�?�og�:���C��M�)k��m�|��	�1vťY4�⭔TQ�C�{�fc]�n����L�li��f���hh#�^K�X�0	Ȗ�gd��-6]F'W����j��F/)�r���'�p̮ ��c�oh?�pĲ��8F7���iI�䯫H�xh����jF ؅�u����)d���:����� ۹̔�D$o�۟�6�ŕlPo�Lۘ^��Ե�m=&����^��i%�u�z��g(Y����e�R%d��]<�g����o�*U$�#�xq��7(c����Ot�0���Sٲ��	"�C39I]�o]�ƹn��$����˞�y���DH�>ǹ���PZ)���\(�5��TN�a�q���i�#�͌��#�Bu���n:J�p�AN��#a�@{:a#��CP}+tnP-&����H���2UY�/���ِc��|y�X	�L6"��2�����B����BS}��\��s���8_�����\A�̼j���ȡ��'T��&[?����"�j���Qmz�6{r�ԁ�Y� W��J2�ǔ60PS�fc��Y�꿕���
.`�k�J��rf3H;�Z'2��/�����o2�|�3�������L��0�MҺ���^y���'����W�)RB������N�ͻ�:x�3������5����g�KyJ����o�M�W��=T�d��2�֓0Q�m��M��Ys�H���P�v�eL-�W�?���!�X1A`d(�$�G�-]���92\`��zYz�>�fe��-x��D^ԃys�mؿ�����*�^������f�����T���[[=^B��e�,늯i{x����IaNy�Ҽ���8Ed���2����M��(�%ɼǮ{(���$h[z���<����J��E�{%􉦤���S�r#�>���Qr��D��*�e+�T���L6�<�w���udw�x�oz�<Jc�U��9�����O��Fn�a_�,'|t�n�Ep6 �}�Lz�N�᱑Xt���p{�%�{��߶������P�&���H�w������(8�����a�0��h��f�`�N��@��`H���L�<&)%�� @�$|_L��o�L7��?�7�9�X�߮�f�Z�z��|9$���?�FqOФ<���!1���
�,S,c~el��n}�Z�HP&�s~ Q�K��#���@��3� '�XrcJ�~TT���^�N��;�mB�J��Y��\L0a��LW4����8��B�K)4��[eH���ʽ1_j����w��Mn�{S%�WOʛ��S�S�����W��쭪��0ۮ�id-�M^rۦ��x�GMs��mݢ�j�׼��If�0if�����KU
����k1��SC���U��z+�-	$��h�mG=��F�l��͑Sʵ�>�q���U@�&^f���?�m��u����r�����Y:ۥ�c����3ߘ!�d��퇦�`�X�j�d�	t$:���7��7&������8����4�Y��=m�P�v�\�;~x����#�Hx.x+�UiG�:Of��p���gL�״���D 
��<&g0�a/]c�O�_@ d�ڜ���7D���[K6�I!���3��Ec��;��nH'�,o֎}2	|9 cα��	�����+Y�]��Y�2u��\'U24s�H�����hU��{����y�v��X��mL�4��lfy�m�&�}n����jO-�B�a�][ t�l_PL��W�L�E���WYh��U���*����z��<�3{s���m߉�f��xJ�0T��e��86.m5����@"��DGh���$���@l��{�0?�:��Qn�Ur�'�e"�=a�il(�j����m�y��{�?zBk`�%�fd�fc�:I���t�#N�;�:Jut�y���9%4S���j�����i����a�*�eՊ"�_�9���З
�$t�H�Ϭ�����(��Lf`	��NU#��t'�����F�*�25��~��0
	I� �+��'�����4>M�C]�8���<�����x��,�*�($��a\����Uz�е�� 6�ֽL(���哊�����U��o��*��L]��b�)N ������E��}[�T>N���j���޽�H(-�է*����,�3���v�[:�:�}������.�04Ҳ_���F�#���!YJ��=�x�L�c�q���x�3B-�\���se:�n��w��\�E4R�/c���o>j��/��4��e�E�܍��/���u�z��s9`�=.�-�kVSL_R^��Q:����lj�WԆ�U��o:AV��/7i��2�ʘЪ�/|CVjůs�b���f�%��EVR�6.%ӧK���` ���2m(֙r�m>O�"��.���O�mh�^Zh���,��g��ܩΰ=f�'�v�sO:C����2?���Ͳ���a-q�Y~w��;�ȁo?_�݄����8Z�-"����eT?0ٯ5��W�aw.��W��sK�WHa�.Z���ާ��_k���l��f��`��";;�@�W^���>b��~xl��/��o���ͭ�e��.q�O���sMH�9��z���ø��4b8T�O`D�ϩ���b�߅�dn��4��\n�ڧ?I�_�f��Z#����&�4\�(���I�B�%�q�n����l�/�;�$h4A�y��K�(��O���/��G�>�Z{��7�g.�`]���$a9㕡p����,������[X��x1�*��%K�SRg&�3H�M�u�a�ʔ��z�[2��vM�T�g߷�z�@@�{�ȀC�=�gx.�����SXV�V����ٷ?�z/�F�Q�}"�X(�p}]:ps
2Z��t�����$�h��<Ɍ �8�aQ;VB�����n�'�O�����s�}F �'m)�&�E&u$���up�6V�V0��̂����L*����O�H<Oh+ltN;��v��	��r����& 99$�{��b.�{ �|����#]��$>���p�)�?�(����}ߐ�n.fv��i��x�a0���/�.�?�`�[!nԕ'd��}o������w7�N���5j ���pmـs �Pjş1P�$,e���t˛{�5h��/�̹.�nݤK�E0:��]@� ��8ϭ{$t���R���F���#P���YM�ȣ4G��g�eH��=������V������֫��=�.[�܂�N Y�X�p0�Ȣ�ŝ}702��h��T[�95q���H}��[���>�&��_�����q=�C�óp�qɗ�r4�
��!���4���~.�W�[�)R��U[�L^�/����6���a��
�ݾb�A,v�*^*nd��#l��H��S�}͔��Lz}ݤS��_�:#Y�s����#i�rJ,v�Jȯ�j��.6�b�	�	Ѯ���ˑ��!��O(8����J#���RP������aՃ�cqu��M9{a�n7%�pZ���	!qӴhO+�4��x$<��}5�{��/73�R8�h{x_NX�5�������&g�"`��eB��1c[������O ��6X[	�.�9}Cur/:��n�ǒV�5+���"&��3��FQ���UoL�Ps���#ϼ4�$ڕ�Mb�f�l�a	1>C{[��^�۸���~�0����4b%�U��u��J����Z�$r�s^���x���r�oU��ߌK4G~���%�choO��1/���1��y(�Mp��6�ޏ��#�ۻ��
譲��ee���w>>������a��u����怢G2}=�HC��}9�,�*�;n����<�`�G��Ė��j�8��ӥR�¦��&Hݖ�y�G���t���a&^oY���c���0�X::^�/��;������p�)���v�#�1`Dڌ����I�a�2:��Cɾ�CQ7�9GSf��}�4�a��!�����g����Y��1�[�+f�����72�i��;�<��|�\%5�R�/&b$ac�3��J���=�vyEwi��ђ!�Try60=č!3ޙ�R�(�c�=9H_���V1v �X��ى�ڏs���z?+hL7re]�rݧ^I:g��Q��>�m0P���Z������;&;ͷ���2�O��(�g�0
��[�X����`���
��˭�0���	;2�E^�{��m*��v�b%i�%�H��0P��oP�=��Uv/�Zl]�)����S Z��$��|�u��=�%�v�j�J����e�m?%x~���Zn`�|�n��q�ʸ�>�����b���^�U��PG��X�����o���=%���g��!�I��0����Y�ق��)��pٶ*N�;�
�� ��O8$�	�t_�R�!�9��pA���S����Sz�O�Ռ�v�藉�򷅏�S���2��0j"�ơƵ 5Y���]�a����A[[�d���k}���S{���0�VI6�5�����$�ڡJ�1�X1s�ή�9��8�������٩7��|�'��|y��E���ۖYg�t��f����c���U��#�72^�����3[� �2�����%��\�R�i���v�Ok�����U��*0~�E*�|�xf9�Wq+fP�n�5'�#t$P>������0%w�j����E�IWٳUTn����+)ǂ�u�ڲ3�0U�t�d?����-��t!�ȡ�������߷��V�eh~���y�*m^�KD;�����s�!w�]���w7#}�� ������x{[W���Ͱx����;<�σ��]�y�����������ʑAŉ�}'���\R���������׉J<���*��qH�~��`z�������g9{�Z9���%<�ʈ�U&~��7g/ۦ��}�'��#���ac>Ȭ+H�V�O:j�$fa����1�:��"��_�����'��)�U��[�h����H����AH�^��!�KZ:��j��P�/�&el�I�N���[*��E��>&�-�Ǐ�&z;��ڕR�ُ�^y,#y��[�}zvL�¼�yV�NG���L ���k`�V�B��FZ��	���b���`��|�6i�F\ʕ�vd�����?c�,�MW����UD|�R�zs�Y4�찶#f�1��@�]�%H�!�E���F�Ww&k���	kl���2�|캢�Ĥ�Y�(�������+{�{����~	B��
zíiM��g��gⵏ�������M�,j}��T��O��:Mcˇ��Ѩa��}=f�����Ҩ#�����q�A -���Y*�wm�r����0�#|V�a�1�������Ѱ��z�3�_W�Mv~�|g�=n��z׆X������;g�@��i�	����\]����)�י��R����w����xd���a~3��ui���:����5�#@�oB�����X�-E��f`�:D\�"�L�.�R����s�,���U�^�"���z+Ō�ҿnN?������/�0�M��ݐ�)p�:�1��cw |�]G�`�T+"����Έ�W۲���Mm~�n'>׬].ϕ�/��]뵧�*�svE��2"-�f`��7��=eʂ������)�O��.Ҿ:ė	�P�Q���������X6���L�YB��+�n�?{��K�ڭ�s �M�����~�\+�d����0~Ѫ)�� ��?�r�\���{�4=��N�x4���F@mw�X��$ڶV��d����8��A�ځe�t���x�ӂ����#�;I)�L\�N�6|�B�^2�E�/��	>�l�E��4�Fb�L�p�)|�Ȧ�x�jf�m�6w�+�\u��#!��U�Iiq�"%�9�S-}��z�?���]��w��0R��ׅ�WI�	�zb9噏d�9���%�EN�e�B����=\?y@ �V^�-�1]��<��
�Ue�tY�x��_�;���.�#D������4��9,�9���Ve@�|HN�3�[场!{�ũ��&��%zM���m�0����['�c-=�(�5Q8��_�Pva�wϾB�&���^��ʣ�x�; ��� !j�Ah��~�m�S	G�9
�o��o0��YZ���1�����O!L�!��>Tq��H/Ĩ/����������j��N����~���/�m�
�����%o��!jj`��F(O^˯,h��R��+M�ʄ�[��=�p�#���qI�@���P�sh���x�dO�Qmz`v��>�u�[IIܱ��;��/����	*�*�m ��D�E�ڋ��|�_�n&��S?m1�S�?�8�!��Uf�����L�	n݅<.{+�#��m���C3�����*��(�zQ����LAZ|�<��ſ"Ǵ7`�k����A��;#�|>�DxAB�Q#^	���o�� 6��tI+���RF�;�u�}c���c���T�In��c�3��kG���$7������.'<Е�"~9�_����d�oY��=^y}i#��|��S��h����
��ݏ;�$ĸƺ��=8��:�lٝ[��m��b��3ԧAg����R�㕼iw3�6�t�3�ص7a�Į�����̦�!=e9i�j�����Ih8����5a���M�fW�7��?0U2�ȇg��v��;[�G���<@ ���/��S0�<{VTn ��"�]1����	��bƯn�/�P�J�S�Ն�Gh&xC�H"��$�UAi~�j����	�2�ڞc�~��+�'���]I~ݱX�YE��a���]д�">r6y��I9�16��Ӈ��C���ﵮ��U!ya_�z��,�%��|�Aʂ�v�T���r�Q(�^u��X�����u�R����{_����x&������3�;�ј�������� �YF<�i�s����������u���&K��;w��Oy��M#���(���p簐��z�!�l_�P�Z����#��=��������w�~�=���Lr�9��wkr�mϱ�:��g�,�5v�kPͬ�}zx��ɩ�P��x  ҡ>6N;ж(gf��H�W���J���0�!�ow`�E���{Kxε�rz�kk5���\7]�{T��n<� ���eD�Wu�X���`�
����"��M��69����g� ��s仳&�RT;u���1^�]7Js������iN�ijڥz\�mi\���s�Mh��[7�x��y�!G4+k �g�>&z���i�����e%NJ�$�Խ�ci�ԝ�<5݇'1����l�0$���K]�p�L��U�����ߣ\\z�2�QS�->�LCؗ-?e*yȹ��@��QBE��w+Q�Ŏ3#�2��Y⣘tW�yU3�&�ȹu
D��w��d�Ha���&����4t�}^%y��P���� �N�׃5���ť��]�2�5�)�d���� -������L�>[X��b����N��:�
�]z]��4�����p��Ywy�ݍ�f����:��A%k�2��Y���0-����@6�]�x�ϩr�f?_A���a��2�l�t@ N�눎-t�Qr52�o��s�.c#B�|\�	��7ih��1⩽ �	Ϻn}�����qWl��˶���ļ�~����U6
�����<aL��K�ͮR���O2>�(��B�k�۟�YkT�G���,�X���;6��?���G��0j�hi�M.�b�-���oW��]�⠿���Cv._Y+�.8�5	�V[��R1v�l5�P��	u�{�ˉ�_QY�Cv��#I�Inu���R���o,SjI����㺧lC�0FME��%UV��֮Le<�e������Y'���d�i���w�	�]Hkg;�d��L���
C�M-9U.�
�q�d�:�_�c%�N��]))��־������,w95�ՓP;�e#����M�0@���6~�Ձ�i�0C���+�.�~����+͑�U��.+Xd�b��,"��$��y)�.GT������Xu� 3���(���S�/Go�h�Ŗ�o���/HN�������t��-����t:.��J�4{م��퉻aG�V��"���fvN��>�M輖rr���!a����6p����u�6�N�w`!p��#>��wo���2����?t4�-V�ru��ߛڎ�@M_��L0�8� jo�W-�},H��'�N���R�v�VM��r4%����4�}�H��
8��.�eBBUXw����o�g�YpU�49-1�4T~�Tˌ-�����i��*�z��p���נ#:-��@�'.�a]�K�눮�]E�T��}��24������u'�}�m�w�>��<;E�۩.^��-����2�^���AX��SS�$-��1��oc݌m�kl0���u+K��0�-����qGU�*=���=��+<-ߺ��4&��û�������W�
�c�
I�|l'����, �vͺ��i��cM��[���$9���_���^�,9Zk�Y��rsQ�u?q�^�ϛ��{'5�5ȱ�iI?��n�~X��`A׋�r��=d>v�����-��n�Wy�9�e�E�N��Sx9��ס ���CW��1�O�v2��{��}�N#�*�x �W�+�7�N��n=�Q6Y�	�%�-��b:ص|�^;l�EH��W�|�JҢ��Y���%����d�Lޔ p��b��Ӳ�O	�l��K.m���F�)3L����V����͈�;���u-��1d����Z��%��(ǧ�V�[��$2O�˒�F-~%:�^�ul���9𑷎@�2���~^(P�U���]S$ ���i�D�R���6{�"��8'�qx/�Ώ"�x(�9�,��K�/+�N�=�>�|��Xt���3�r���_�0l�y�Zg�5��G�z7.骺r�W���XiV�d��41�:��N����|���x��B5O��LO����6�SA.�}�u�@O7���5;ո�tm�-�s���?��/R�����s���Ɵ�8����F��?Է���R��<{I���<��[�̺A��8(S�b$����Ѣ'�`Ց��"���J6�cp@����}�@ֱK&��ۡ`BXk���U��g��~���6��{WC�^K�z,x����[���S;�_1
�>L����\��ŵ���a#��d����;PN�C�t���`�����?A=
����[ӌքӠ��i˛llnS��m��>�o]~W����Rו/&�����Bt�g#	�.�X��X	��*�Դ��*M-�+UE�n�:���2Rƀ��K1$5cJ����l���m���ߟ�֤e��vv?�3� �X��@�ؤ�흗֢���P��[�B�PՂ������ kM>�m�.�S��a�����SQ�}�p�1��sۏ��\a�r��_VcM�������Ԓ=d�ܡX7����@��M��q���� ��N���2۫�"֌�W�أ��v�Q��]<֣�E������Ҳ&N�)T��,�"e�h�Y�=��M���3��
9�����tK}ar��]q|�8���ff��1Tl�{��UU���Ř�T��#_�S<����0O��Ͽ�����zL��{ON-�<�F�D�r����+�)�pu�.���q�AW�	C�^���]�!)�����e���If�<K3���<\$���K��*W�٬�3��8��8�K��P���m�2��.�8�����۽�ox�N���l�9� r�}�~���cL/qtf�Ϩ��(j�K�$�)W�II��,W�kj����AW4��+�Qh@�o�kR{���T���uǍ]U�c_��c�[M<8n���4�]�ښ�/���DNO��eco}D�x��%md���ٷ�b5Z��-���sL����c��fh�ڧ��,�=)W�,���~�&�aQ�75Ot_��o975Fw�@L��e�j���g�U�!�QO�k$�F¦ΈJf��&	�ӡE���@�S��^V%}�iQ]�ː���F�;��G��C����Ko
�I@�o�nl��q�k��/֯��[R�"��	��051=	�`���'��/p���]�����gV�|�bY��5睾]F�}UW�R�.��D��R�
-�tg���l�q�g�.@OL`oB_�6x��c��>���� P���;���k�TAo�į�>U��!�'��x5����@���?r�}&6M�kk��C�h��mW��l�?�.��%EY�T��!y�x��漘�|+2���Z�|"�œ��J�< ��w���<}����ՓL}ƹ���P�?�������*&D�Fa��4��׫���ɧA|�$�&��b��p�O�	�jЕ(Ǳ�9)*b(Uz��|�P)�U�c}��<�pt����կ{����~�"�¯y��=
����Lme�r��Ǖ��Ё����Yh/m�&,�UGN�����`VYx�누~1b�z]�&�kc�*����)ۦZ%X��߿�%�	����?�[ܟd�����`�|�+�;���4Z�$�u������$�6l� �B���39��J�B!���9`.*>EM����L��@)k$��*�բ2�n�Ƴ�an�(�2Tz�C7倫�<������7�gh�W���-����?q/7U.�o��43&�Y[n�	
z*�����^oK��sQ$�h�V��N��yV#�v\��k}�2ď"��.� -GF�p�6�����|ܞ�h�ڀ����'xыy��=���ǣR�����0f�^��bE���3τ_w���[5Yp��l0�v�>�	�V��p%e	3�7GEwϏqN�8<�+�y�<(���0ߌT�3����F��gC6�v�?�ڙ"�CW�+\� gL\��ɤ������Tk��e>�}
4#S�~8-�+k���*�nyU� ��0)�-��2}\@)u1E�y���l��G��N��R�-�0��Q&��`����q���܎d�% r��gı�'�.4�X��ʟ[����Bi��r�b�w�3��1y,�!	p�Unw��+��^��3�@�5o�<[)���i��+�2��U;�6"��,���
�i�:��x�[�Dw����( ���A�U�h�>Q�#;� �S�y֚�����	�X�V�z�r�'яlν�7FWyلS�둖wC�<�=/�S�;�yו��a0�RN�Y�׵[�aI�|�nd���R ��~$?\��̖lk��b��QJh��FQCn�B�1֯�� t���5���+���������Yg�K�<Tp�����^�9��e(8=Rء���[X-��,�O�t&�3�g�<�/���j��|��s�v8�h����A��	��|���u��Iw�T� 
��ߋ&����[�\:�����h����2Y�l3�^��uS���(>��H��犥���������擷u�������B��J���-�"�Hk��!oc����nu=\b	�7^��6t)���TV��C��[4����|.��hd=�l�AO�`��>����1���{�~�m�
+[��ɱ���oC�j7��t� 4�c�<,�2�����^FqByO3��)�h�\cC�lɣ�J�xk�nd�x�BO�}p��V�K��w|��	0�/s�i���驅�\c�u���wf��hJ�ȓ+�g�hgy�^�bP��a^a;9�I}<��ly�sS�s rp{詺Œq>�iVE��/ �O!9z��',I����G>S��m�п�P��ҭ��c�]T�$���k'e��٠n�Y:�ٹX���}^�������8�<���]2�7����Rl*-���B��!��mD�"S┘�{ ��f�2�t#dj�gr���zR�F�Kǆ6n�ٷ=_[d���.>�+bG���X�Ш�;�(}<��4��h��h�:j�5��J@�\�����pSdV�����m˜F�9� ��=�Q�N<ϗ�	;�t�K�R���fI�E��A��J���Yy�C�;Kz��I͙ F#��mEo�v"�TR�0l��mlA��E�)�1Va_�|Km/���+hC�Oj)_�F+��� ny(Z�$��F4Y�'�{ms8C8C
]�VI6���R�R���:A
�$�5�llՒ�'V)��W�(@��<Wr$2*6���OL�>t������Sb��h��t�*ͼK㉠~��GP���(��֝�d���S4V�򥓵NF�1�0�*}/����q4��ZW
�:z�I\@N�;�H0����3�:��-?��g����S��N¸�/wd^�0;޹y���W�Y���<���g缼�5�&WЩ<�}����ޗ/�Q�|@A���C{G�xLw���L|k��_��l����s�g����S|$P����|�E�N������5�=��L����E��sĆR�K@�?1y���[
�>V=W����νĻ��������D��������j���r��t���I1�{}uoN��kOH�]:Y�ct$��T��o�@���B�,�c2~&6��┩��b�+D�,֍�>�D'����XA��o�^a��fk0,��z�;KA�cE���u���~���x��Fq�*��P���Ơ���x�s4S__�O�[m�?�Ĝ�­�����G��^�[��tgl�[[�[c��j�MK?-[R]�ʣ��~o0�������K���15nV\lMK-�tl�@�b��:��7hy8#BO�l���g�(�33~��O��Qz�B���K��'cg����f��b迟J7D=����,1�9TX�0ձ܌����ԬZxm�����Р?�j
��brN��ko�VZ������m������߃"/co��E�����w��� �^�#+%�{�T4�h�<�[W)��[����Q�Jܧ2�_>�;e����p�=U?i|�ǁ�:(����Vu�?RU�j�sv����/��_{<"�~��J����%���q}�������-t|çc'WBRwJܺb_q�P�#s��<Q%�D��T-�l�t�q�����l�r*��vj�������SSh�]ש]Z����d��V6�y�"ҘIue���N�u;S2�������H��8^x�=^�����ӾӜ�����/n����'f��wݰ���`6۟o+��&fW"��)i��#v(��d�LGu���u�j!��OA�F!�Ϗ��e���<F������_i:[�iK��I���E�˺Z
F���MW���oy($��1kV��Y�g������]�c�C�T݈0�mX]yw�����Qq�������9tmg1��p�?Xl,E��,��N5vw��l���ngD�4c(Ɋ������RFJ�@��Ul��٤h�z�y��T}�5-�4D�[�[��l(�i��u�ː�ُ�[�f�V���S���FY�n�0������}�q�%��oU�-㤷��U+����o�O���ӗ��y6�$�/�`F)�|٠)��3���<qy�8���'�wY���g����� _��w�+�Dݹ���ir�"��H��x?`�7��n]����qj��\������m��k4��s��\�?n9GD�I�����p�\�*��:Yr#�y2>"��C�H�N��f��:;���VZI�b��n��15P�C�*"�T�~�\��_$�� �7~��Z����sV�29|��**��}�ߎ��!>/��ӉVҌ�v��3�0��	�¿�?���b�ġ�u1h\�J@��En� �u]������m�Z�=�I<NÊf�%���?��Ǡ�fs�Xؕ��Y��������33.i��-F�
KJ6L��ڮq�I�J3��J��hV�7<v��dx��+��5֎�wr0�8|%��2L���6�㡗s]AN\�X9���6��qe�a�6+�t�������UC�E���_�{�\����|�V��{Zr�)�����%d�s��"���Qa����"z�Ȫ�>����OK��S����n?p��.'��u��cۓW���E�o�fJ�j~�#��7����F��qz��q4�� 3%k��Y׭g���u�����{ߺ�14G��"�����kǍ�'xm����Cw��\�j�  �[	\��ɡ���/י2Dؖ<W"g��m��?XlLOx�LC%��p�|���4�iM�"���Up�P�}N�5`ZF�|����;�!&>Z���U/pH�������g��^ѩؘ���AY���+��t �;ў�{�'�U}<q]��=�� ؐ/ �""�5��S࠰\���Cj��G����?�K;2F#��ݚ��P�dR
v����Y(���o�a�T��5����GT��wu���ॣs|+-{d&b?�����^���f�+ѩv'�wДrS�{'��
�b��\îT�iz1��p0HU�'EI�$'������m񴡹�U�>\؞ ����	��x�d��J����Ri�ѩ��Oc�O���E%��-�M3Y�b^+�$2Lk�?~̌� ]�V��b�meC"�k�2�KN�q�Cx�랛�qN����QmKA������Ӄ��ڭ˲r�&��U(���,0�,rL�����mװ
1�z!�x]��V2x���Ȅ������ޓ���z����H�rJ�a;t��n�vl�\�ro��BH
��q�+��^Shr�\��Ƭ���Ʉ%��DxTĠ����.��Y����<Y���L��l�)�l;I��r�����ˠ��<7���ʺ�M2w����T�bh'����s��:�!	�z�F3���J�%����5%_�^�$l�&�t[�2F��g+���;Y�/���(P۾Yp����T��Et˫	�rb�DOZ��S ��7���^~��^�;�izK����utio��]����X!;(��a�e%8�րփ��2�C$;��)���!�'�7o����Z����@݉G]�כ�ȶ��V[��_[Y���V�A�<��k�7=�|�֪mQC�x�౲��K�T}�:|�οǨ�CWW��q����+e(���F�x��m���b�Ƚ�Gy�
u�!kl��w� ����T���;K�v�d}��)
��7��>{B¼�����)��O3��K��1���\k��g(i��rr~�ؽc��+G�I�j�[��nB�ֺG�y�����Y����D� *�siқ�*�tAzG��Ф(*R�Ҥ�t��B	��R�	=��z�����sfwg�yfgv�eG�`<O����-��j4��nJ�Ns�����*��T�j}�������9L�_�#l�� *��Қ�y���+i���o^�J�m&<�����u�*K�}'lYR�hD���/9�W0��ĕ���;���3ʨ=�7Or|4��ݔ�"}V� �:��U�o��oH;��>��𫴠.�?UAfǚ���WM�C�)��� ��Ld��c�P������80,� �P d���t/�N>t�ғ*U����},����O�����;%+�5���2����j�#S�/֨j�4���[b1�#�n#Jf'��r��>B΍�k?��X?����f�>'D�=����g�&�wk�u���)�Wϒ��qT@M�|#�PR}[:��y)Oq����R��������$��H�*�f�Dd��ùyav��@��Ã���石���=�(��D��a���#E'��ς��H��Y+�-��*ׯߘ/Pl~�QKh�]]��P��<�C�����V�S�y?d\y�͗.w><����d�]_AG;�p�I93sY�z�����s��Ʒ2�iR�j�VpBf�i�5a���5���숷6|��o��F:��a#�M|ذ�F6<:4��f�����({���ѱE����a���K��c�!g��~p޼׹UYi�|��.J"ۗ�W������G+�cR�����@h���{�Qe��+�^�#5K7�-=��Y�w��h0���}rٍ>�Wq�H����X	�``��ηL�Z&E���bX�hi��/�������hb�4<x�<m������}z1�a٪�����ui��e�[��w-g�NR�*�m�E+�H5I��,�T�byA%��t<�������%Ӕ�?��7Y��Z�ĳU?s3���$D��%�{���5�~ �3;{��׫��V�Za_�$����_��L�f�O���oNg@���Ѵ��2�Q�R��5����Ρɣ+��2�`]�����
���G�O�l�D�7�z��ƥ��~�U,����E�*�:�o�_�L��t?G�n�?U�+r�l������z��4/%vY�����s4]o�[��l�NÅ���Q,ᒕ�kC�T�2�kmk{۲j�����]��?���d??xb�ݴ;�N!�,>�z��=%E�]7���_S�Ôb۶��	�2IK]�u�G��긒�����z:���7�Դ�S�4;����H�Ȟ��}$�U�6��<��֧:��GX�ۧ�d��؂v聨���TI�w~���K���[�xW�^�����@`�hHkr��[�Q�%�,�)p	.�v��[�0ƥ=�pH�����#6J�ŝ�w��v]�V�{ɻ-�����b<E]aӓ�L|��(q��m^
��&�RqU���y[ĭb�ڭk���g:����Yi���\Ӟ���z���7��K�?�PrEyziD!i�KH���*�[�$��́�R�8F'�z��}m�S�Xk}��#'3+*�Dt��ܷ���)b\v��7	 z�@�l�n������rqss�g�`;B�u'n���T)v�W�Zz���Э�/� ѢT��S��Ҧ+��kSv�xF��J�8ϖO:{N_5:�η�
�>��y�靾���_z��bpe��.��� ����z݉��ҦVL��ұx����!b��>�z��v�.�(t���B�L����Mn��ó��o�	�42�T�B�m�As���<j�%.�T<ؗR.�!�um31~��>jFEl*V�KqF% /��NoQP���2��
�nB%�z���.;Nq��F���~݅�����n�'��h�+ :�,:a�٦����1`íg<$ưj���=�7�p�;l�\T�p>��Pq}\��[¤?kY��*�@��,�o b憭Fb���ɓ�	��;cKx0�3���n��u,k�VvU�$!鰠'~>6,Q�����ס:���j���{�y��U UT��#�&�-�|�AyE5~BP�Uvm�N��x�r�tH��i^�L�D��5��{a��q׮�}�bK%m����Kx7����m�0F�͎�}&5Φ�!g���V\9R~K��T@�9�i�{��e:�&��3�U�){>8�cX�g�huY�9����B��z���Y�9��������5Ȱ(!y�_6��մ���n��V���K�X�>N�樛;��R͙�͉B_�#��c^�^�Go�k�A�;HB(?�q��1�=�l,���ߗU��ouY}iL�?��9yRt"�2��D���g���E�����vu��ss{���^�_���ւ@�RD�B� =)�Vy���vNq�����9����TY�@�X�7��SU��鍑�O�X�Տ��������aʭ��1��h43�,�Q����c���No��7?���c?�T����M9F�4�#!�;,���Y62X�,x��.�>�ʟM���s��T���Im�YVْe~j(5�O��>����A��'�d\�c�բ\d�|����l�'��EY�\�hU�C��1bgS�Mw���Iw"��k؆��:`�&�����P�i��R&=ۊ��?��jv|ѭ)b� 8/���|�l2�JB2�RW���ȩ��>�J�����0�����x�Ƒ���[_�G���eZ�p[ƌՋ��ݖM3��Α�Cݏ�I"c(s!����{�ɨm�>�$�9��E���>����;>Z 7`'�1l.��.˗ݜÛ9ۛ�%ҁ�9��l�>i����w�
>�5Q1O����혲���PLy�yk�y�`vTO�H��Sx���O��0�����~W�PW��R��zBᓒ|�,�prh���r�A=�K8����h�!e<Q�C�c.ĂApd(b�5���seK5�!��J��S�r�uN�vr��"`��ڦCvF�W�D�hS�M>ԧ=�a{�`Sݍ-�.��"����v�1u2����a�����O�L疎C8!�l���k��P��YKk�e�x{�pꪢYٮ��Li����O)*�}���N�_��˲�r�fP��n}����o?
X���t��q|r���}�����1�^���w�)���>�᳔�yQ�R��RT�ҿ�SK���:��KY@ �n�͊����M���=�����n-��U��v]w|Ѿ�׾硾�X��u������݊q|}����Ψ
�x��\���-��zOL�K�;����5�Jfk��.���^"(k��*��꒶���]^>Na�E�-[c�on��sky�*u��P.�jse����St�ѥ��m��u�%�����N�U��ELwV2�M�YYU����p�� *�����EG�����-��9g��[`]{��B'q@�DS�Q�<��lڜ+�u��=�a� }IL�������'�=��^�����2o���lU������!�G `e��4��sO�k<8Y� ��]����/��2��in�Y~7�kr�N,��W�{���Yo���doz>�`[,�9z�.���eO
�$�����tVj�VU]m��k��Z�N+@a�k�V���;��O|�_���/?���l�qL�~x�B�Qh�+ptV��р�P2G�f\�W�2w7R!"+�3��<|�]^t���6~������.��NG��F�Ǚ�>� ��u����s�-^�(�(W�~<�n�k��i���3���(J�.�;�rrr�,>β24����(�	�嬮��y�bTB��j���0����������3�>�z�(�Զ];�'ث���4����h>|�l�Ԏ-��5�j~1Ea��'E��9��~�{>l�ܿ����*��!F\�yx���k�T�}r!�aAa�ʭo�t8Ek�ԉW��^;-�/�{ZY5���f}�$Թ�ˎ�zk�<$���Ѿ@*�`̤�57{�~t�kr���V5�YmN��j�l��M��w�A���5��ٻ��\ۻJ�I��<1
�$o�A�'�6	�%��˹/�9��N���H航�EB���-r�����/W�5!ZxrO�"4'��wO����	sc��Ө��fZ����e�1���5���:ӻ�M��C'H(��~.��LԨ,BU}�M"I9�1׫C����G̗�*A�f)��0�+Þm�w�\��YJ��( 姞��+U֫dޣ���p������Z�c�� �O ���$���lp��Sྜྷ���R'db��7�ˊ�S��yO���� <H{�h�sf7�Y����]���>X
F���#���o��R��~�l����� � ���*��V��N��hi� ��i1�{'a��RQ2�Q��X��
M���Vmt���W$�q�	33��䥥F�Uwd�.����y������w��b=#�B<�*_窄�=$c����,�y�{�B'n��J����$I�����%љ���.��d�ƠÕ�e?����FP�qy�vq�)oA�j����fm�����!夊C�� ��='� ��2�w���`��0E�c�U2�º�"Z!.�-�E�R�f��6����� ���Q�"[�ں���מ�iz��J�8�\i��Vl�y~������1����s��f�y����ϱ2-|���)T�L��P9�s���&��<���%Ĕ��%��Be�0�,�m4�� �u��S'�iv�y���r��׶X*��1���v���z4֙ARg�p��%/���S���.k���?\��
����ٳfjߴΨܡ^��Z��pX�*�1x���fU��v�K1>	<c�mKqԈ-m��E����@�>�	�pp�\Gf$�{��f�U��ʇ\ZBn���h��j�W:�O��z4jMc��a9�9���'� �� 0�tMה%|��s '�9�鴜c��#��F��Ƕ%�����J|�B{6i���NK|v����������V i8��*���[j��7-����s�/=U��mVO �l~���T�6д��[��P�U2�I9G1ʩ'AǏ���S,�����*���}��Ad�=��Z��.f^�B�檲\$�z)Y�[�fh��v7���^f����o�ӯ��Mwǳ�F������.��K�Lgx�n�M!���p��Ś��*x�'�,�zVB�AQ�oIC��R��K��pM;���t�>��Q8�u���C�s%��CԴ�$i'v-b8W�R~�tMs`�񂝔�z*��(�jl<
)�����JK�\�qt��s��g����E�pr�8>�P����.�7�?�~��/����^%��?�{iy�YK����p�F�H�4��r<���Ղ�ssl�S�ƽ���va��i�2������r�}��֪1�x�s�5��:��MJ�Sy����
�0l�\d���	�����ܡ�][A��V������ A��>�Y�\�u��;���|l�k����4iʐ�d>.|�]	��c����\Q�2|W�!z�c!��N�����;g?椖4b�B#LpBWߴR���ͤ�F"����j{���N`d �9l��憻Cc��b�LG�l 
6�v4�\��$��45�S�АRŴ�y�D*��9?���~��ڍ��9�T��ܖ�CkhȒ���}��K���{�q���<���Ӳ��Mj�h�����[3��>���]i7�{l���Y�������謞���~�)ķG��g�����7�x�:�޾�\��+�?~ejz�E���;�>��-V� �]����,'�|��7�0le�01��ͫ!�(�9O�n��I�z�j3��첲]��SC�O[�|R�&�����9��I���G��vV�!*o�V|SȺ��tù�⮪�mn]�~R���g���:Ɉ���\$�依�.����;���f�õ���d�G��/��7�>6��!0���B�w}޴�X<�V����*G?�{/�tY���U�2kNqUp�
�3R�Af [�����?�ꖲ��l;i���n�sE^�^$�=,z�8TV���r�Ǵ�&�\�J�R4)�lV�h+�n��ģ���	8)�RXB��9�9^-b��6�VP�Q.S��-!޺��Rg��흉��,��%��v�����kb��4<� ںS[j����?��<'���%��O-��2�9�<ļR��h���
oib5Ϗ��AY�]lT���Mp�p�$�M��>�ʉj*]քjЄn�T[hu�pxD{�Dg���l�)I�����5`j�j�a�Ok|�u[ ��*���a����Y\��I\w��s���Q!�,��:Z��������)Ǫ�]�wo����'��j~V븁Zk��FM"���T<^@X$��h���� ���_���%t�s]�]m��C�`����n�S'J�ةj��0Q��Y/�,?9�Qag��NzfI�?T"Q)�p��=�v�iDYѓY��mfn�}��T3��Sz@��յ���k��ʯ/�J<�r|XP��R�X�ϛ�I�x�M�aa�u�wy��_�<�ܚpF9q#�f5�%�bH���Jq��W��u�/ܿ�0f�͜Q��r>&:��{�4����X�՝X����F�P�ڮPR���oz_M��Rr���p>�T��_Կͭ�{�E}i���e0�Å4������3�c����������|X��+C�D�Q����딿�S�M�����߱ۺ�_Z\D'(F�-�c1�z�?f�L$/sO,[��v�:�E6V�h����F��_GgȐ�p��x����2hL|�f	&)T�u&�zퟺ �74�Ң��Uq�S&���92275�c۟��7�f'��IJհ�o=f�Z�oY��ϽKo�����Y���3=<��C���f��s��MWgX����AϜ�Ծ����]���F�Yr���b�
IhM�v�8��A֜��8��>�c���O���|䪝Ɋ��覱����l�*aR�U¤II"}Q�,W` OIy�,�֪B�j�`�FKʉ� �Uδ��}��M��1iF�~���pa�Q
sw��"��Qh���KX�"���i�ԹF�f�3�nQ3�6�x�d�c|�SÃP�6C+�����=���6�c�#w�/�B"���JWe��Z��K��
"���JRx)�e����7!��nN��֏jw�K����4ȗ*�Εk�V��W�#�ϸ����ڒt��"���b��z��W���?[y�=���3ؼ݇���)M� ��ҏ�/,���o&����OA[Х�S�ک�z#k��a��Ψ�`�|bХJ�Ԭ<s��o��J�jX�(r������ Ί�o=A�(ppD�<Y}Mԓ|Y�"ohK��^&�JK����TŹf;����l�Q��O��d���m��^8����,x�?��"#��hv5�\���Y����#n5�h/��X\U�-n���Uy&��I྾�T}"����#�Q��&���[��
%�C�Dai5#`�a�n8����^�e0��b�cf�~6�6�W�Kֳ�ݟ
�A�]��� ْ��!*���9���E�n�}d�} #��pĲJ�$���pvl���`NR�
���䁒�3)�n��S�j �p�9�����b�)&�v���4c�n�q�m|�����b8;�i���A�4㖉��d��������kۜ+3��>��=n�:�DӺ�A���������C3�
r�2�E���������j��`����������7Eu�d>А�(\�E�����e#�$�IhH1fv����ؐð�cͽ��<���K�N2#W�kNDre�!v��aTB"EM�Rw�Ϫ��a�F�HO��ʆ��#Gg=:�	5 �s������&...���/���˹����r��m�5&>&��J��ǬW;=ˌy=y������\�2=Ǵ��ʄ�{�.���*9�.)��X�P�q�~K"R���L٩��.�����iT��j���2�Fiu��g.7�����U�\˯��q��I_��xz
y�R��ARS��z�\j���q�u�ӃJ�(�W�G��&}퇾~�e0��L�My8�{�ҊUoX���;�購s�D%`��E��V�S�nk�r
@>��˪�~tK�=:�MM����뻥 �s�7��E���X0L��V���^�|��@̩��Xi	����8\d}	5iM{/#��p3}�5^!�c����\O�����a��?J�sa�M�/6J���[�qL���[���4��|wt�q.%e/&��O*u���1����jI$�q������<�;(;/� �2%e3_ |M���C:Iyi��7�3��С�Y�{�%pL~�4�7��0�w���6��L���,y��W��޹���xB��i�/(��$��i�a�n��NT	J�ZfS�k�$rX�ߐ|��cb��h>��~�Q Iy��^�����|�c�0��ӝoZ�q!CE �r��Z����GT��D�N��X��]��g��l0�t���$�df��vQ�\tr$��|Va+��x
\�}�+j�;-@��2Rh:�!�Y� �O��YT��]嚝��� �Å|����?K��~FC=���f����32��`����n�~��<C���le�H_O�@�S�7�~�Z����1��f���u6�zKa�4�笽fN����	@��������Z���fF83�n��!���!e��ɮ����;���o~��z?Pp�-��%�R-"yFr�ΚhZU��tg��Ә7��5n!1H�uXk?4L�B�hi���0u��
qy�!�^b�4��P�F���3&�r��{S%���B�ڰÝM�3�١�a��^���{��J�^n
�;T��9��R�w����u�������Q}�)�"n���J���/
]@3���w�m��<���U����L�y�^�?��y]{��H)�~0iw�ҪR�k�����ۯi��L�,ў6�"�g��2^���]��q��n�c?��4�
���p��Ui�G&r[	��w@�x�P �H���	���ů`5�v��YK` 2���ų�ſ���b�����7/[
���s�o�L!%�d��Q�S��#��!�w�/�ϓNRW�%L�mw��+'S��8u+�>Rݓ[P'ڶ�-_�浂�DiO�}yG�T��ˎ^?�{�@;��ƶ|s翉k�]b�|�y�ͼP�X��S��]���e��� \%���n�J�=��nTV��MQ��rJM=Բ*�B7deRQ�V�-���_���R�� ��9\/X���U�i�"������e�u�g�A# Ws��[�nX�D�/�`���1`�����ü� �d xN7-��n� ��|����I~ ����P��%#�*{�)d�G"^S�Qx�_��SK3�R4����!���Ct�֣K���Q���G��8���߷��-t��N/�6n�d��L>����L�=K{���u��=�L6m��A�E�����������<����FTI�ګ�������w�m{�����焑�7���@N C���355S7��i8w !�~�v
>�KL뗪���~Q���PTI�ٳ�{�>K�T#���N�.?N�l�h����d�� ��~�"b�e�Ƅ٤�DY��^�|��E���ZF�1=��UqP��YK�N�������O�����Ю�n��x����m�~�k�B�r{e\_;�Qf8�n�O14�2H�'�Win�$#f-����Ҝl����w(j�mml�����Fl��m�3Y:L|�&-}��(�X�#��=kR~�u�Sܗ�t&>��F�߾���>b7���%�K��M��\��s�w�N���a嬞�M9�^�|ز���K-�qz����o(pwc"i5�B����kLhGD���u:ڀ�"̐P�_��#v�oG}���ϮUP��r236��-q��}�NJ��u5z{{��o&>��]~~}��ݽe]��<� �YX��74 z�պ)�%�a$Ǉ�t\k�-��*�$���hj+�O�Ty�����xi��,(h1�͛7�����b�0���l��]�8#�F3�=F�K�S-���30�:X�En@����NP8�B	�?�oĈD�E�7��T"F��~&މ��X�c�\v���V�ͼ�`L҈�J�y�g+R�PC@=V궝!��e�M��A0q��syu�`nn�1���2�@U�B��ᨴ�u���e���V�V|�V?��P�-~�/����2Ѳ�x���-k����`�1<=;�ɱ8nP��'z`��ѽ�~x���I�=�jYI��Yj�n�55z�_L��iab�Y��r�/�sUۃguM�����-OzO� w˓�V4^����x��\1
9q0����8�OǮ5	�iɚ�G�����W4��ġ���?�5��������o�2��!1�*#
=��M�	ֺˢ��1[*�{2!0L9n�%)R�C��t|��ma'��hή���m��Aһ��"��Z�}((I_���zf|莘pFB���XڊyE�5}`a�E��r���M���Kx��""6�%ޕ�x�B���b�ҮV����Az(f�%~ �h��<�PAn5���k���*�N���\2
\����x��̐.������ґ��Y撈8�m��+�5B�'�,��)�~V�7О�3�b��~���i�h֐�i�C���$�{���=6�pة�_����ͱ���+��'���>J.|p�3��}����^r?�A�!�t�Ŀ ͑h����2�Q���'���e���`��o��mF��x}�k�������	^.#����Jt�^S��ؤO��O�;x�2.رtFJ��؂�.G@��q*/;�F�"x�%Ρ�����Gǵ>��b�����nt5h���Jܒ�,��xAU̜~$��JLb"�,����|U�X-w�5BhtܨÙ p�d��]$~g\ Ɉ���)	�C�ʾ�\B����H~��󾽭�{�c!�
`�{`^�,���]K���siNui�Rg���A}$;��a˛��΍'�����2$��5_%��i�A���#NyGt���Tњ�)%��I{�k����P��5Γ�� �p�L�+5Өp�^ml�i�-�;�t�s��E_l���ZqY�\S��Y��hcs�/UF�n���z7���\|��!E3�>����kC�m�(��>ND�6n.��П�M����Z�Sꀵ��r��<��O���Cd�=	�;�c��K�a��H���r`�iOѡ���[�<�/s���/�+|K�r14}[+��1�|0�g�v�7b��Y�=�v�����ȅ��s��e��b\k��u.��C��Y1����Z髹��l"�^싍;���V��g��)Y!�:�.��d|��S���wˠ��`��`�-�ϧ��W̆�_�8h�ͮ�� ���Nss#t[��xqГ�&�B��T��03L�]�Q�J���Єrw�}(�'�<��;1��˂�(<9Ҥ�c�/��9�B_Y�0��r*�ɭ��*��ݗ��!:��s2����둠���Y�-ғ�(�g+��Y��~'���ۮ�$�J���ذ06���2��%]Km�U/�G��o����Q`a����V�_�>PQ\kX��u�zd�������zD�}�������ԧ���K�=]�H@E2��~�^:�3�#Ӕ-��2�2�Rq'��NصR�Jאb:>
ǯ��VmD��Eٞz�/����@��u�T}�2Z��<�9�I�!uY�k�"�����q^��]�ao��O�B��Rz��)yH)�K���wy�r�_��8dj��=D>hf��N^ÔD�U�����>�~	L2%���s����:���;]%�'�jd�֖��t��x�Ζ~<�&Y�9%z<�J�M�Τ��!$���d�o�ʴ��b��^�KW�0ĩ�ax�n��=��f�lx�%���j�w��bV��_��.Sz��!�BS���<5�F�5���pRKwZ��S�Ub7��v��6������@�w2���@�c6�TJ�����lT�5S�&93DMl�l�|��GK��b	!6U1���
���ZZ��W¯W�����*�.���� �!�x����u�(��H�/CWZ�(W\
���CI��u���ᥧ���\.�̀�w��Mk`�0Os��~���z	c��rL�eS����R�4�f��;6���Bm��Ho>Ar�j�|ᯰlxߥN�M~O)����| 敇T��ț'!�\p�oci������%�t*�RB�w� �`�����%�Mڎ�t�%�bF: ����U�j3�{�y󕳾e�d��
��gN�(S����>���v�2Ȅ��G �u����t�Tڧ�Ŧ���.ױ���9e���g�ݾ�<�?�3_\)ͳ5(��"� 1F��V�(��6�cE���.�(d������磋�-�os�[��>�F7mG�ӎ�\��xE
ڹ�������M�&]-jŊ8����c(���z�^�j��w�K�`�o����K�-+1�R|����"ي���BQ�f��>�ޏ���F�w)I��`Bٖ�'���sp?���:�{��������۠�̌���L��mxOD��y����w�홻ܾg'��� 7o�QF.�/4U��m�8�ke��+��*(�Sb�����PB�'�����'�����`����@iH2��X(��6y�$�+��\=ՔP��e����g��:�d�!��ә����iҍ!����Y;-��3�����Z©�2��+^�ؿ�i��䢖 ����W�n	�3%�a�j�].������dg��n�N�gδ�4Six�6�>5�#���x����s�;��2��^�p�_���6���ڙ���Y�}$nD<��_H�.�حu7�k���$�s�.T;�ԣ5�%��\ �uh�� �,��o.�2�'���+_+]/r�X�6�&��ڧ��i�����I�׵�D}��R�bHy^-|����	Q��X�Xڭ�~B����X&�q����o\^����RD{�G�uȏ]���5�dƅk�1�լ9�}�SY�Ӻ��u����ag�
�����=��/�L�Ǔ�}�9a���WA��5Ͳ7|մ;�T�><q<��$��XO�ц�[��"��O��$+�-e
��G�-U�["V�,.��ޤPP!Y��5�V�1~o5Qegqَ�1���<� l�_#����H�W�%`�A�z�Y���_o��ƺ�<g�a�&�ي�.���3_���RI�8A-��!��Dq|Tƻ�Y�`)=��}faI�ߙ�v P���vB�����s }]�	hZ��ʹY��f�j2��`�B'�ʵ=WL���
T�gnr����ߠ%�U
�e_Vb���?�-�+ɣ�����LYu4Z̿�%��(���us���V�+!>�3x�]�;��K�=A)�LƤ�]�zlG*w<�u{r���<s�)��_5�+=�֞'6�e$�#���=���?y���֋�8� |k�~O�wT��o�4��ٱ.m�"�)U���(����ӗ����o�H�x�(,=Z���)~]��䦫���Q�4���b�Dbym���y)�9]D@�hג��%����F�ۍ�B[C'*r[	�S!Rq����c�OW�??s����`��B㘼c��µQM�YQL���ѳ,���~>i�D��K��A}t���oW�Qk�l	[R͋Wב���U�q�7���>4�蘮��}�M�w�V�KPFt���U���B�%��lFO��OcO��8�Z�?� �R����0�1�	d4I&<	����ݳ����7�$�('�d��@0�Z%!��
԰�L?�=��d��}�+�MYkz5�dGt8�C3OR��[�T���"�
M��:y⾇7L���:��E�oڤ��W�Z�����>����W�F�|���-�zH���O��!k�c��%�=I�<���7����y�����6;��SX�*���#�G=�~P��1��$n���^q�&$�`� �[�Vڰ�=�z��z�QCb�2��]�if�
����ů�%YT�ǜ,R�r�3��C/��ܖ&��OOY�0*x���RO��Ӗ�/m긴�����������x�L߼��sHu�v!�*�W
�7btO��Ti�F���$�-�AFk��G��xG�/����&�T�9v.:YBbQ>d�{j���i��[&�'��_ ;��{��z��]��&�{�Z0p&a���H��!�"���v.�<���hB����s�#]�9;��T'%��t�'����$�Jj  ���F�GL-K>�i51�2��6Sȃ�k3x������B�>��v�	����� ���rn/[�����L��\)qR$7�䓩�D�h��0���7��m)��k��T����6��vG���$�ѷ�6Jȓ�h�����~|�X�9�:���G��[�g��"�M92Rԃ;�6t�}����C%jūwI J��{���}��ߡZ���s�����){��D��V�V��a¹�|��b� E9�Y��]�ƥŮ�Ƿ��M��߉,���yTn�kP�h���iBV�!{�>��Q���+wEVY�8��O4�n�U��e�0ԑޥ�ea�@��J�ӂ����_m'>�)�J��1ɑ���A��p��WO�8�-ʻ5�AK�A�R5�u0���1�5r�0Dymz�W��4z$f��]RP���u��d�q`�JY�l� (z�\����PqE��)�\�����G��=`ex{R���/�����>�n�Zfj*)2�<� YN��</��S2N�ͱ���W:Ը@Ɩh�p?�4�a�z�ljE�sk�38��.l�FE7F�`�Ɍ�w����$wPP��KO{\	Xb�;m�MQ &3�a�2wyfҾ������qO�-����K?���+,..~vws��Ц�5�[t3|K+D���<�S\F�'��کVx�ފ���y3෧�
�L���� z�㋔?�^1�!�J��V#
�1�"��#���6�������G1�콃���V��WC3���f�N��=�O��1����[��\��'�d��W�ƻ,�XV��?� �]#�복�A�Q�Ϛ*̷ӽ�7f��|��^�pb��?�@��G��%���{�G�'�-�.�,d�K�)�nn������:�fƭ��Vj���4�'�ԏ4�A�O֤5j$��en���2r#>%W�}���؇N�, ����*��B���w<�^P�@=4m��'�NKL�����/�aT�z�`�>apsI��y/s�*<�j����.�O��`��+�C�^��7<����u"Иˠ��L s��G��3���!MZ�ɯh�J���,�<�*�X��� ��r�?�Ey!��كV����=�	뭿F�X�g�G�?�/w�1Ag�o�l�Z�=M���ڢ�k�Ι��Co��HЩ�&�-����C_H�ǳ�9i���#�-p��%��H���|E�(����[�Q=7�<q�U����Qӗ
T-���N�X<�����s�APT
��1����N��.[#΃d#�F���g٬y�*�ލ�@$�x�K�\^���@㫂��}��J������mB�yUٱ�n�v 8&9����ž��A]��CG���$)"A��ˠſ�+�KB�"s��߻�����z��+d�Q?yQ��//fB3�Nd����̸O�$�W��`s���E~�V_�!B�O
��h����W�����n��R������7I=��H���<~���c'a����ϑ����K������v�.��P4e)qhoC?V��W�Y���S0��sbڊ����74�Ɏݗ���f;d4�"Ϋ��"�T�d�h	�+��%+KP��N)��c�+�w1�N�K��d+�V������jħ�S��f�]�z��������]�����,����p�z�-2��v��9`$Z��z4�V��Y�l�XG�c�J78�n5���˧Rξ��H�4Ѭ�c�uQ����A�b�`'���(�ju�����b*O����%����v�L��7]=�Ѵ�&`��\&(+�Elz?6x���p+z�U:��D�����;�z�)hc�ʶ��	q`FэL4����緻������ЁM{G�N631��#����0:>F��D���?�Ԉ�Fª��%��LݡJ-$�)��L���t7XY\���\�ď�jYBg�lЅL(�NT��r�@1�<�6��O�"�b
�=Q��Ή�5L���Z՚S�s�������M�k�N�X�^	l_�/NP�@Ǻ�;J �H���f�d0����ŕ���p��G8�w�b� ��)8K��D ̀V�((-�|����aVZᎪ�W=�Ƌ�⒫^��S)W� ��r�7������-pJ��"I����mb�خ:�V�}���jR���[�^?? L$�c���WG�u2�|�=/Lv�'�=�n������%k�$��%|k'���G$��IY�S5q��S��Q���b�{�D!/
(����xv+�.�I	h��%�f���~��
ı�����z��$%%S�C.F��N�2�����]�5�=Q��8�ZLm\ɷ��4�,s!�2�o�k	�YГ��(yt܈�[�WxV2�?0�'?��2�*��"5�@Ww������g�7��$%��{	�^9�����-69T����{�M۸��=ѩ������2א,�6AӇ��#EA��"��@|䍗2˳����=�}����F�傖���-���������A�o�����@(KZ����$���#<��4p�5��S�>jbgi����ظ@��э�oPA������팼�2�2��׮�YJ��-t&"rl�44^���⩽�'�8	����{�X.n
S��gWؐl׳��S�_s�ϟA
��O�E�wJ|͖����\J<��FɈB���l��71��n�`�u�W=�kN��^�,v�2kGF�M`zw�m�Q�e����s���Ez�"�2���V8�|�clơ�͐e$�i�={��ܚ�N��2��U<NE�m�t���3���q����J�iF�}n�Z�$ە��������#����\�GSƯq���Ur�(�.n~4q����r�3^��@%��\�l��`�7�j��߻P���ε�%)2�K�/������l�ԪCx���\��	{����D��������I���/���<����x�{Pw�epg��[�V>Ʒ݂B�!'��3s�T_k�y�Eׄ�bV�Y@���( 9A���d�%.�("y���d�9��9�%Ò֕�d�����u�Wu�n���N����	�}�~�O�$�=r�����x�Ҕ��ft��*�k�"�eW\�G�̩`�f4�J1�7tw�a���Ǆx��Α���G0�����R��@P��}���;<�X�~$z�1�&"!��L��S7xJxm({],��տ�ӛi0�M�.6��⡉Mװ �*�[d�w�+�BbS�Ӓ�gn��;��a떝x��E�spE6��{mY�.evt+��"�7Q>�IOz.�y�	Z��,��j����� ��7�.ގ���~D#`�	��'��l�g��M߿k�s�s�.����\i����pS5�	6M���6���n����ޓ��PZ� e�F���F���a�<��*���J1�4E�)�4=�GR5��� ��e^�;�z0^���sm!� "�(ȟS������:��¯I�¥�鄧�>Q��pU&�>�'���WO��V��\�:~(.ؙ���:�b#�{��-��9�Q)�S���{)�){3]���Y���=�r�G/u�U��R[��2=F�+[���g�j�}9�[���;��.�X/�f���1�}��qSƯ*[_�@Mt ���,�Ԩ�#����"�C�L�|Z*d����Jjt~��X?e3���Щ[`0�.W�Y�+�U�*6k��+�S3����Jo�+����>�3
�sJ(j�F2���x�2�c�#��X�Ձ/���H;��M�~n��Y��JY�}���is9N�3p3/�,�(��*�[�ٰ�<�z�Lg�kw���j^ax��5���H�?��P0#+,l���*�NM�:pu>��`��?-O�=o2�6q�7��G�!�\슆*Q�z �x4���'\�0Sc�'���
U�,^�Dc���VO`w���P2 &z��R~� _-DS�!B�'A"�W��	+b1�_j�է��?��ٛ�q���Т�ZVqX��S��6'���2��M�ccn�?i�ۧ��AM�j��ħ�v�"�Tܣ����vHv�0�݊�k0��wvx_r�WK!�W[�����Mp�*�˫��Ɠ�I���Q�������6���I���l��°t����	H7Q�u_ �8���w���|�]�$���8�r�oZ�g�ۀ��N����o�̺���%�!��u�a}P�!�糒t��026[�)����� �MK�/@F4 V�~�<Q���Q!�V�9*_E���������X������D�Q�ԉc�"�r|�h�06\C�������U�{\>�'�4<?��e�e��y-.�t��vɼ�����cw�v�q�Ӽ���8v��(̱L�>d�����!a��['��	�GZ(�m�� �i�S\dN�_w���zab#Ya�u8�P����9��7t���򲗷��ϯ&"�vw�����ѣ�5���7�M+jY��;�,2��m��*k,.�@^�rz�~���
N���8�?���ΫwT��H'0�o\�R��R��v���0zM�>������$�/����~{�/����h"!~�"�(�WSH�*t���%�#�3�h�
Fg^��F%�RP���d
7��}�?|G](,0�|�0U�BS��C��sJdT��2_u4R[��f+O�L�}rh�A9 ́��Ő�8�_d#��48�7�և4�8ع�����7���"o��w�|�.�ݛ�ƚ������"���t��0X�0a��:���J\�Ũ����a|��iy� �I����G`���m�RCo��v�j��E~$��8{��r���-k�� rA^+���i��>>�I��(CC7�1vc�N�]��.�*���M�w>~u&��+�'Z��/��;i���&0tMS#�n~�����ȡ�
��E�A���sۑ������7.�C\�I7`���k�+��3,>~��iW����>k�-q�ڞ���|���tT������]�*�d�kb����R[�OG��ۍ�}��1�ؚ�,�,'-`��ǅ���"�4���s}��󷎀�lҎ?]<��2�d���E�	������=�۫uFU���
sիBS� K%э���SS2xxGZ����S��"Q�f寢<����h�����:�]px#�=�H�9�"��ý8 �c"UX���I���26���4�ֽY�	�P�������s��.e�BL~r�>�h�� �i����6�E��EIir���&�Ws��R�st�\q0z�N*�A�{���B�
^&s����k�����ˡޑS�ԙ;�{5�t7��J�ILzXw(Ԥ�Cq�
a0�����4)��j{0�X~=�1�,�$j��7����tv�T#��xC*WLHK��;t�5&��s��;�y��Z��FP'�4o�m���
J���K�\�E����Nc��;=�{�:����dV�_��Vqm�C�i�BF�Zr��2ׅ�P0���?LOۯ����l'�$�Rt��x�����63�#�J�\ʝ�a�
�e�^l�n	��JZ5v:_X�Ha�aTecg����[�RYZZ�x{�~¦�a�_x�X�3Q����D*?�����?����睕Ŭk�ϊW���?bZb��P[�jAex�r4�nzKe���DڳC3�ti�<�4���q�
��)[�C���:�J�IE?RTT���5�/]OU��i����g�;�oJ��n�|#'�$��" 7RCu�]�v��B���:�ұ��>V��ͯ�����g�/̽#Q�'�\���^lU2���G_�G}Ԛ%��ZV�LY�?�NVڏ��g���N]��f�XP�e۸����O���5��=5���pS��=Kt~Z2�"��*�	�ި���ƶmIxp��H�,ahX:CC>��J�I�ǂt��m���ɬYB�EKK�@���+ ����fV1�*��1i�1�$�S��E���{��t�n�m6�J}_;��k�+��2�I�-�@�}!�Y�^�h�:�[�1��l���q��V�i�Ga;���y�w`Մ�'9�b1��O�����|խ�5����S3��h���/��s/���	5.,��xی[K]�iR���(��	�
���q�vl��;�i&Q�Cg�pO��6\x�Zp5'}�O��y0��J.`����V�I���v�^a���?��m����^��VOs)�60��6W�����V��wkG�0E�\^��2%	�+
·U�'�h�ђ����j�G$�h'�z��Ɔ|�\����"}�$��V���y�C<�����$����ES�'��<~�ћˉ�*���^�%��ޠ3C,p�'�ٔR����Bo�د��!�����u��?>_��eP�7�9#��T>W�'v��!�vUJ��1�o��?6ے!�&����񊊊���Id#�.����C�w�V�C�Aܵl݂���Z�R�����^Vc$���
{���d͇%�v%�봉	���{�%|a
;��*��mhb�Y⟟�FL���lm�$�"���tF������ݢ�I��g�<0-a*uo;+�>���:����"���Jg6�����Z�$����9��)�]F��-�������^��9L�~̮c��e1�5�<��ƀŶ}���DB<Z^6"�?�`�b[�JQ�&˚�����������mC\9�!�I��A)��i��9����s�������ih��u
�L�FN�{;E0:�ִN��NcHm�����R�/0W�-ˡ,;ѓ����%�=�����QF���_�����ؔ� �'�illf��7j&Ō������'Хk���l��F��֓!�{����]��[ڸ�M������<��AZ�:G�F��5����o�::1�v�J������ڒ&q��w�[��� S?%@��Z��Kd�M�B8L� J	�����Hb�������b?�\F*�Z�<=lxm����m�����KZ9��|������f/L�\vH�:R�7�X�
��Ѿ[�1�..�!;�x����e.e��H!:�"���e�im�Q\c[=�^]�D���*�o��,̗Ŕ#LCf�(��bOh��u޴e0�a�����o_��a'�ǔ�zޣw[�Hߦ�1�l��ʔoMUJ���T�����-����,p'�D��N0r*,({	br���A� ��%KY��焓�����s�!K�|ç�\�.v|���n�F�i7�~�A" �����r|ٯ>*��p��\���<F��u�|\T[�4�,���q�U6h�X�	cr����^p��FR#�nJX@C�˹d�-{4����c`����f�ذ�o�.��s����e ����l�6���Ad?n��"E$Jj��NH|�/�=(�`7��*�i���o��!q�l���T���oE���#��|�ǹ�c�����a���ߏ��:d�u5����������J����%{v�-_IdX!S���q��j.�j�Tvs�Qo�#�?T�%�Z����Yh@^Z`+�Eo�l-��6�ڎU�B���p��	��a9�HP��)n��H���]V.�.g����9텭�N�2L��Π�����-��}���c숙v,),��u�;��n��0��꟞��m?hTa���$�8�m�#�����b`�(��ȨQܨ��T?�@��۹yN&�{�2-���]��:'q�#�q:��?�=�tU��?�|X��Ӽ�l�X�q4��!�>��3>��׫�@QjC����f;�%b����_8�j�^�̬�e��/���.G���g?�(���?|��<
?�q{���z?&�÷Z���F �5�,��)pL�����x���{t���2ҹ\�LW[1C�ȋ�;?����' i���;��d[S���%�~��c��M���X����xkiO�qu�����S�)q��Ŗ���{ƍ"��s�{_)?@Hk�~�1o��x+٪.�n�Vh,�Փ~Ч��#j�7����L:/5� R�+��OIt���A+���$�rlQ055u�E��Tc��}�( ��_';�Y���}�~FZc?�&��C�J5��(K�2��GDQ�d������QCy:�!Ӕ)G����'kD�]�G�h�T���)������%m�������۩l2(����\������"�}� cV{	�,���5wQ���|#�����7�U�)�d��e2>b��\Ú���5wQ�z#ƨ�Sz�q�K#q�?ck�	.�Z{r��^Q��k��8-���r5�Y�|������������VE����gpp|�n[s�ɀkrڨ���R _NS���/�%���I�1�ľ/�/j|I�,1�\�H[�����f��h9�' Cv���qE��2�������ҿ��S���)"�&)��A��/V�61$:���m��"N-ʂ�}m��ā����7c4�/&U�m9��G�#� 7n��Z�?����Vz����xZ W}��ɐ�o��ɏޝuUZ�0p��|���Ǔ Jxh��O����Q}�����ܿ��R/)���^��^�?�\	Xr�*�*�B:�c���y`q�+C��{�<�p��;@w�́�8=x8���E_�<fr�N��� ?Vr��[�6p2���<�N�8zs��#7���0T2��(�����~�$-�	.�-��Zs��i���i�M�	�_�0������� PlI}��@�\��[�Ec2Tk�O���eT/����¹ԝ� �xVh���G��;��k����镾t�'ڪ_<�cK�1� o�h��덎`B� .4m�g̭�?.jq���6�EzS�	���_��M�L���q齀�x��~�@�\j���@��o(�>@.⵿��0�34N��<~]]�Z�6Y��'-�=���L�3*kW���)V<95�Mf�) <�w$�����?]k�5�!�ބ�<tӗ m�к�K��|sY�@�6��×/�Ӱ׸?��Ou����Ī=:���V�7#��A}������o�����sU�W�޼|�/��� ���/���_=���~#��� j����+eT1D@h���u#�.��1�0nbdj�ym7n��|ݛfF�c�&0���z�F��l9Q��Pe�2.�eD�<���<�f�>���w{�̓䬬��, Ȩ�.R���#�ςՆ��Bt�U^	 �pLQ:Z����H4���{y�eja�������_��wY�	��	J��0c�v�C~6������R:g��H'9u�Q����d��K��퐅�=���I�Ӳt1��~��Ν~<PY�����Q�M8�.z�~̐갴�nA�F�{r�~�b`��!;��Կi�lLXv�����b9�d����զ�Eng(�>
�(���2���ڿ�K+����)��Z�N�G~��h���I��O9�x�U��Nw�t���������7��Vݫ���sqY���n��k�R|�,[�N���������� w�}S���	�e?���g~N��j�Z�����-����7	�UH��JC�m�xU�á�5��#�[�X�J����m"d��̜�*ಈ�%l�<T��CLM��^-X�x�[^R셱7���
ڰ�d�x��[�س�<��\��g>n����L[�N��3�ul�.2���T6"]�`���F�L[3�ZQHN��{hX���K�k��R��2�T�|_��aAV'�N)��[��z����B�[� e��rr�[@�p@���s|,�M�l�[�����}�
�_$F)e\�W� ȩl9Ri]�r�� ��4��;r�R��k���5[��U�, ]o	��pv]ɓ��{h<l���xs�
���k��ﭭ�"�ׄh���J��V�����72;�^�.7.�2a��p���*�!���3��c%�
��;�G����������Q-{EO��Gl8.h%3�Ķ4�]���V�Y�!!���r�f�͍��~9ݷ��u�1M ��Ӹ�w}xm�ˁ��pU��w�oŜ%d�Vlo4Q��¹O)��crԢ�1��m��z@�'��a���,:vںe�^���IF��l�13w`�s�HG�l��lJ���f$��A�Ս�rާ!�:��j�qqa�k���dh.�&��p(urྡྷ��m��z��&��×�r��v���39��&$�*���o��SDJܢuP�3]���oT��j�Q��;�rr�`�K,&�^�-.!���LC�I8o�|����-���4��T��,��n͐�<8����~ź�3�y_��`��Q��bئe���Y��+6~;k�!��|����4o��	���L-�p8�~���T��R_x\�)��>.��������է��A=�����5���� ����āҀ����d�u�{QVtV�x�Wj^�i_�">Db� �,z���-?���`G���x�*�>�b$�V����[�tI̀�[���ߵo?�	�6��{��M�ϻ�{�u�g0%�LLr����ڊvS�~S5�����;�l��ֵC'ר1�أ��⑩���v�#s�ɛ#�s$�������,L�K�Y����<ƚ�a�MBF���W���"��O�۩��c�xj�<�ڙƑr�:��� Ԩ��r�I�ML?�%��Pf� ���@��B(AL�vM@tF�; ���o����(��7��:<n8�)lMĚ�ƅ۽\�J�А��z���<g.0�����Y�Q�㝼�{Alz�N !�@�[�ɐ>���T�MU�E���DG�&��M:{�"N����x D�>�ˤ�.�dV�oe���׭h\{:]g�m�\�\����(��#�ʈ��6�z�̜�y�7{���=��XY�F�+�ָe�k����\w���\M�Z+@��ե�Z`��r�z��)W���8.9�fk��P�?w�uX<�fXBi������c�rU���}�i8$��l�9 �[���ߣ�r'%Ŕ=�j��=s�H�8�����%x�x\�^2�\�03�@Ţ�mw���pi��̡��q��);䃻
*�_�<���m�V�Gƀ!C(G�i�yK%CPK#�C��f����H���i�ӑ���>�8H󢀋tZ�h[�x����Jm�.���V���|�_C����b�� %��D�-���InKq����;��f?���`�EvR4$�k���UU�)Ǔ��YX����2!��'f���-D�t5?6-��R��mR����;���2�h�DeZ�gw :Ů#Њ\��pE����x�9��[���d\�H��)�Z���p���)Ba�8Y����j#dZ�p�^kw��Z��`��4E�{�(;�VB�]yK�M?z�'��Q���~lh�b4?B<�P���C(�?t�iU��x0\��d�y:f?���/��D��Q웒��03��|�MH!�'���1I+Ї^S�(����B�5rU�C(���-� w����Y���3�mv?��~e ������P�pKʷ�������r����r�7�����o���5T\��Jr�]��I�O�����m��>�� ܽ/g��T�j
8�^��-/iy��j0Gݾ�=��,�00��f��k$,w�|�2f??3[��_F����� >����?{�1���Qf�w��k�/aT&��5�Snb��c*fN��A��J�Yb�NFJ�&[���|�ѪɎX��K
��r��Bh=-W�~i�δ��M!���਌e
;6�/�e�1�N�?JCb"�'K�`�Į8����V&�ݙ�j=�?E��>WZ�!���SLb�<��7¨:����(�V�Z���Ab��T��-q��RJ��6~����-�1�M���OBYᲦ�� H�t����L?�_�o	�gYt搪�
��`@���،y\��x� +&D2A��T�U���r)�u�1y��qO��ϳR:cM�8��C
,��b:�jnt��W�~���� �is%��>5O��ܨ}t&�?(!�"FVm���m~�cUJ�J�2���	
�L����7g67V��N8y��9b��"P��o���V�f{�Ӧ���k�,�.]��':5��J�c�v6k�����g�x+GN23i���d�ƴ%�5��d��L����{��� *h���{�@?�)���<��B?h%k���or�����o��:n2������ ��k���)��H�r0g!�	��t��n�z$p&��GL\�L$�mح>�xD*L��Q��{���j��g"T��X�8�Rۼٟ��������|�H\�IU�zy}�E ��?����M	ߛ?�M2��.~�`��<�ޑZ���a&g�pc�'��I��~�Y�V�Ч��"˕��q�𸌘%�\��W=W״��JgHUn�@�M@s==�s��%�sM�� `:��9�Kp�@?a
�<9e�)� 7*���(X̏�����t^0}d���葶a����� q�ޝ�k	��
g�k�7kFk���A�Y%�t%��OKm�A�Q�-�����/����,�����Гـ�K'��O�l � �aV��cI|u+koh~�/t��h�k�ޛ��k������'�<��+����������L�yr BZr��(u���+5��k��T�N$�_�0>q9XI�'՗�
����-daӃc�Z"g<� ު(��9�N}%0�V 9#73ZH��Ҍ��1�^nJ�� @�~��n��P�O����A1�ǂ�@ ��&3��
�y����A�����-�KG6�@�N������9�~�ge?�sFGz�?�x��c�Rӌ��v�zy��n��}-��j<Н�'�4��~��Ta�7� �/����P��G�cEu��;W�	���~�v����9�ZȈ7j.�zd��b��QO�.��NZ;���9��L��N�ʷ�����ȉ����y�^Y0q��e:�����V��$`	�-~�@�K˷���#�g�g��i���0ݦ�R��t�>I�?�f��X�)Vp��a\��"��h�`A�Eʟ������zd/f�4�j�N�R�Y+��\l{���m��cK/��	]��`���I��A<���<��H�~u���Rs�`���t��˥s�9���b�=�����g��p�@��n���c�e�'�/�2��q�� �����;C:�t�q#��Ee������%�2#Ζ�@�"ښq)l㓟1���XT)]��.�u�Fyٴ+��b�&���.�i�e����ڷҹ4G�k��O=���MS��7LQS�Ou�_ɮ��P����IP�U�r�$ܙ�+y ��Ps,�+��zx-@&��<��%n�^Ex��W�o�>�.KG���G��#E�A��W�	�2�c8�7b�(�59�^Z4�K��<K�>�@�_��P/��;1�����|�A�4v�q����X�L	x� J��	��r
���GM)_����E���À��B�&�܅����:x�hOw�ݍ��+���t_+���D���K٢8�rM[�!yE�`B�JjFz�������
u}�C�ߵL���m/�"P���1ꊑ���� ܮ�4��2f�BWfޣ�x�����]V�r���d�{�|+J{̺r���ߗ�_42��-�2{�Eѓ����pu�iܥ��(q 㱦�\ZZ�`�)�r���n����G����m�*&&�0�Jd�B8���:��IeR�$�o���M��e��h��a��`c��!X�\	�m��dΖZ�f��6j�a#M+�����U�{x�)C �6?s�N����/%��MJ��Ӧ8�Y���?F}9�xȉt���"���D7��Gi�;�V3���k=)r�b|��u`��ڙ�rǖ-Y��'9��*NV{!�t��޳�dڦ�����׹�O�zN�q�\?�=�K��7�B˺��8p���L��^N���}I��*�p;I�a�s*��߿�`v� ��_�#YNt�;�J��&	��(K9�G~O����s�1ÿ� �=��ca
���x!+����p�M �Q?����S�%��KC�j}x?�qn߄!^Ta����Ҩ���"��x�hڵ[Ĵ��m���v9ۤ���n�w�E���xk�,UY�BR���6ǆ�R���8~�ژ�
�bq\Z��.Xr�%}�t5�:}��Z�E�.���M�Ai5%9
�)E�G��>���P�?@S��#���h�1�='�`��Mӈ�I���).o<A����nP��!��:|����M:�����z�8���V8[��B2uK*я�CTem^ΟF�d*	�P�`t�WMx�]�&�YL�1E��������X� iզ���g���h�P�8n�%��uד�M�*���0)����z��qz+��ȹEm}/k*q:c����J�T<z�XJ5r��%��0ҍ�8[�t��l�_�0c�׫;����-y��7a��Ap-�܊��x�!&��.2f��p����jҊ4y�5�0�$,D�{�5`- 󨜚��3��p��c;�!dk��K I�����8Ep�c�p�Zi~�Բ��Ҵ��� �܅��ɾHq]m�r��;�|H���|/�f�Z���駠qn��i����%rW�}l�Hi��O���k�۰�F���Z���-wO�S��VC���i	���ԡ���·kC��cP=n�l��=51/S��(l'�	�|�ʬ�:h� r��u]�!樐y�=
#�Wk���~�&K
9�%�bF>a���.��\���Κ��y<�aUh�븣�a���[9�l� ��d�Ŝ_(ߠզk1#��`�Π��v.�%�U�
���":+?x.�tc¥��vy���h!;MZ��E��+vW1`x11���X���ǡ�����0!�v������Ǖ������T^�W)�B��EINRy˺�>ek�
4�5y�1sv�S]�d�psSW'�3(�YM+x�sz�4:��ڽC�5��Z���|�'(_A�_�E�Һh����9�	�`����p����?�1���S��?z��������(`��]�]ۆ��S���)���)����@��i�9QFC\f�W؆�Q+�11��ǉ��}���eY���ތ�=���*F��2��c7��s� �]3�G~v)"Q^�X����+C}7Υ��mхY=��d6����<�&ҭEQ·�JF��Pd�8Mب�M;�߳�v�K�H{�I#��1����mi"�%�^������������LL?�ҵ���V�z�����":LL�5�)�+�3ߚn��9A�j���O�<��\�nN���2%j�#��tS������}%���U��=��o�-�镽T�LX�J���)F ��@^>�Ǧ��/��(_?�m��'����B'f�����Hv����E�!�/t��v�44F�P�dٞ�ᯌ����i���������WK��/�������8p�4�X�c%����[�Zց[�Fv��)�v�-�=y�,T�8>�XY8h���Ȼ@M2:�Xa{0%��P��g\�@_�3�u$��$�y�+��Z٥t9�<t��F���d�2�=�e�{�s8"������8n��<�Ȥٿzem��(�����X��Q���wg����$�n�{�݌��x|f�Y���g�]
Nw��تjJ�W�Hp��]�
J�=���9]}�5ٻ���ɡ�P{��ǡj����� @�����#�^���`���+����N%�©�����J�̹Q�/?��&Y	��OE�b��g�D�[�N�X]8���<Ef5�8.㩆<P>s� ����qvjg_�He�oSCb�����N��rv�U����-��=�wm)�~܋�'g��^[�ȹ������3]ݢJq/RITȱ����Z���cgu��d��7wzܴ�S����<�1T���<��7��UO~���<�H�ٖV���z�^z�1q��f������ΰT��a*���{��Y#q������)ߎ�NNÝ	��ߟ�t�ݎ�.��?����1�M�Ԉ���U���bh]�?v�x�\ �߀@�֠ W�Y��O�[���&��n/Sa ,H��`�'�:��5�CC���k#E�!%}�3s�.��0�� �������y?7`��U��,�?ۈ���ٳ8��n �������	�nV��օ�Su�AyPX��������ԛ�s�6G��)lE�;1�*QBʋ�nf%���C>R�����RÒOXE��a��:�W�k��V/Y^��.q޼>ې��ľ�L�3m�Q:4���P*J��߅o6�G�nbS��b��i��[F��V+5-�ui����L��07r�c�Klv��9��m��,�aw�Ku}����^ލ��)�ָ�;�V<��p�תg��{��}�S3�g�Y=�a�'��gɶ�����E�e/:�F����VJ���Hk�"�\���"���� ��=������3������#���u�p�`vZ��W��kׂs����F����{�\Z���:��p���yx�F%��K]�0��d�/��Q2bm;ܤa�	���>��F�%ס���
�΁�� ��آM�4y�A�:VSS��Q����T��ؽյպ
Ov\�Փ"������1�й��f>������[[œ�X6�6٢�<)� 6"�3�ٴ?�����V�f�89�Au�����F��zY�XXۋ94�B˗w�P��ce%�4l�xF���iJ�<h��to9^#��<����ہ�W94�e��>"�Ct�3>�B�J�I��H/�}	$�DJv�������L��=vsw�K��][d������s[bW���N���ﵽ�#������7%%%�#�3Vlll3
�����F��*۱�UvH��*i�GX���y����YI��dQ�bKi
�$�*l/����>�	�$%'g�����v��PPP��nmn�(
�y[P�UZVf��I����b2��u��l�vs��c��D�do?�b��>4��~r�@�=�m��`Ŵ0Xȵ��:���+�g��t��Hi����ZI��_U(�ͫΠ�I{l`MkT��f&�K��R]SW�P4�]]M�c,s;5">�k��:VCŉ-HM���ͭ����������˹/�_r��.���ׁa\\\t=�c��<�q��H*G3�p���]�I`p���@$�n�R�6�mm�|�a��`�ޞ�o��a�f�	���a�u��h}{{P����/_>h�no��	*$�����y�A���n
B�wn}��͢��6*2��I��kT�]�%U�f�ʫ͹�.��r����m��X�}��oii��֖T:~�ߧ�>�JHN^�Rd�ET0��n*+g�u���,SNE���V��k�\{��0]�T66>V�έ\�Bn���j�5�B����F[��ttĤ��j�
xk��TR����]�������Ru���Z-�M���G�ٙ�v�����������.��T�OI�X��䑍��d��==9"����~V�����7x'I�/SS���j�6��	���ώ5�NN�}����d�;z�/22rfbP�z���"�血�lh��s�5+��Rpcƹ��"����P��0�e����;E
��݂�|��W���E�_KJ��\�����Q�����(+)��1��}29&&H�=���p�m?��ji=��OW���>_�#����,[%Y��s���;��������`�P�9i3�r+�lst��Y���iQ�����۞{$��yk~��jc�:��\�H?(((,9��b���{�ވ�4��:�MGw��k��B&Ǆ��~�l}��MW�(4�#�g^R)����rH�js�7��C�;�a�U��[��wChiҤ��KJo���yQ�P��s��ːk���`�/�\UWd�%K#��%�d�7�r*���e
������b�|���3��+�1���s-ѳ_�$	���6�:׻�(��;:M�̰ !%%���OHD/қ�ceeU�y���68�9�&r@.��(`7�f�St-qm��P��C$}�`-DAQ�Ǐ緺��҇������_���<m����Ž���A��=rf6AJ`�z�"�0@qy��5��~,���{���*�(�`�JTG>S�yb�jd(9f�uq99y��X!`����k�d��Pݾ��vUUUյ|gF	�? h�����4�*����Oc�dVj��2��T]��㕍�_f���J+���'=ۚQ��oZX��>���ʲ�#�����kn�^��k��4������bb��6�Th���׋Dmpqq�R�ӧ��8Ptp�E�E�1 �r��p:��TM���Ƽ�����Ҡ�rd[G׷tY�j�c��
��K��z��˫�v�"c���0��I��r�)j��j+�M}�w٪)L����5{��f���Sb>!�W/��5EtM���YRb$�{wc���lw���.yP��5����؛�Ò�*Q=�a 0�����:��w�[ӚN�n�	��ح��?@p$�R
j	"/�����>����q7k��b(��ĢW�.G�S�a95�����(�~Ǽ`1��ᑰ�;�����5��`�4DMf>|ٕl�i�-4�a|r�R�LY��yX�����mÀ���,J��\---��۔'�u1}<
�,Wt��:xȆ��6D���"u����W$�t괣�d��tx��D7�om�k_ƐjbK�����w�^�����$'%�)�b����"䧯$㰍��]OOG� 2�I�7�^]"�쩋$�!N������Q�z/�#BG��?&�f�ڞ�ђk���	g�8��������]���Ha�p�Bg�0�F�xكB%�oCy: P�3Y����ï&P<1#\~˗72c���i3��I�(�q����
G
��
KD����*�A��)��SJy�b,OibXz�ށ[��ì5Jk33�b�����8ͧ�'�+'�����!	��^��9J���%�#�C04���h}�L��0��I��!�E�Ѵ++�ʤF��^�~=���L#0����1�V�mަz(�4
@[�C+���p�Jܧ��E�߿_��9/��B8\�4�J���`ꗮSs_�)2nu��d6X٠�L��p�1WIyr����G�7R�F���#��k#��ce
rwn)���y����Qo��c4�a��8��m����&����v�����6 ��T��Ag�G���w�0��^�x�m���&%������ʹ�ϵwI�#�^��][�,�Z|� �` D V/�}����@�k����K<�v��j�ni��W�z"K;f�?^�<Ν�n��
C���'''��-����]�>�}{�z��if^��حَ蟥�
�{7�̻^���I�R�2��,�/�T\Q�R����U�	��Tii�}��2*x����4��m�j,� �6X	�C��tT�S�qZ�n�峊�,)/oFt%<�l)9����A��-|���yxx��߂^��5k��}�I�w��/"��f��H���L��B������,ʱ9�["$!v�	�߹�ZL���0-u'�C��[o(�=��4�����_���S��[�3:=M��=�_Uh�pO4`���1?:z�n��5��Z����Vo/\?i�S'����NG���)�p�?ڞWwws{�^��X���뻷��BL�����7��*�L���Co��7�D1��!�'eK�-�ifk	��DWٙ��$�l��D�D����y��8�6 I�J���W���;�CR���y�� [�M�ȔC�J��)y]�_�S�����B��~�`�_@�7'�Jx�v����-�r��5f���֣j������~�f��t�ƍ�����G����I�:�}�A�m�^ ���o
ر����4�˄�gb����xw�*e��ѡQ�|�<��}r���l3�I����T'AR�srr�6vs�¬'�^B��c8�F����mmא���و��T+�'�3k���@7V�� 6��&�T]���"��17�ů���y���0�r�y�:\����tr�A����,���x�V��{�Vxd)�!����3�tK<:RVEEE������r�Y&,���ǘƓ��7���=WL�~�%R��'7�[f�HGb� n�����L1��eIDKP��Fv��"$$��|����%M���3������K�Z�_D����k���>;A 6��Ll��2�|+�|<Ip�p���<�^��9�h�%��_\�eTM.H���N�w��$���[p!8��������]��{�7k��:	�i���#U�ϖ?�;��|m���fW���D~�~�***j�FL�g`��rw5;@ŷly���-�Y�a8ג8\�����HX��n��\7��K��78�H���H�W/�ￗ�Rq 0O&&:	z�#��GV±w\2�=���W �ޓhg���;�o?�@���>^��g�t>�nܲ�E:�'�J���V�Բ̓ɚG�_T��J���3ƭJ�����S��IBB(�]�׃~�R���<���X [�XIf��I���`�ciU_=a����+%��ABBڑBJ���\?O���������Fe�e�'�4�|���}W`hq��fKӕ�*�R� ��Q�EPů�_P2��=t����B��>Pw4qwk:��'Q�ݻ�^�\�b��W�ԯ��5��7ǥY���p!4:��U��.@��8YSb�MU��D�r'�{�uL|�T��ؿV����n��'w��Q���6|S�/��xピ�+������M@7;Z��%qZb�K�e��sˡ*����h>�����%�	ei�"r�ͥ�]m��|�=5�|�V*�p:��\V
��x�ʧ/�ru?)98�9����Mr� [z�5zp�������h���,x����[{j8&�w��� ���tz�L��/Q����X�2�l6�0�C�?�QDDFV	
��>�."a ��`�����2Pm8u�ll���kX4�k-���;6�pA0�C���(�Q��K�KK#�h�nе����!�_�k�bA��� ��O�[���b�=p��G��fm6�G8��9����	�~�	Ѿ�k�G�м�^_wg��ys�t:^r��kr� 	�¶�i��ϯt�%-��R�~]�MV��xuON�a	*,�T���|�ϲ�^gAF�t"���y�_�Oy�L����X�Pl�+k�����~W�ԟv��*D������uM���P��K�75�)B����:���.����^�Xkv�ŭ�
�v�hs9_�s$���F��پ�\�)��K*�g݇�o���.�na�"xz� B�=C޿��iƥ��)������C.�h��d�X��x��J^����aN� ��E&V���Ɍ5��Ӿ'/��	�}X��?���,G�m�����:�� �O�T6���_�j�2R���FXJF�D ,:E����A	K�e�n�"G�.Z(�Z�k �Ob�W����K��IW�Wu%@QY��I���)BMP�B��qu//����O��s����G^Y�&i��U���0!��g����5�&ʀP�H�c��_U;E���+�M���'����W;\/+t�tX����� ��y���vQF���B��n�/�;���Sz�&�Ro��jR����Q]��v�xv%�s�H���d�D���*��Ko�k��P�$��EdI	�~��^����*���aI/��ƚ�Bur���#W#�[���w�8���T-~"����������:Ý�����x�T��G���{1>x�s�p[[RR��(�U��N�;��I|{C���'�%��ѓ�)�����kɧ->�=
C��`:ŋ�hDçx�,l�nL��'�fNo�!V�L�l���[�������O�j;d'ҕ^��a`a�1�S�[�㲘���_pLv(0�����)���ƫ�$2�eetu6���h�Q|����MMZ�+���z:>A4��TMn
JbK_}��V�(��$�N�R��P�rf�SG7����F�EP0z�s��\���LI�R����)]#W�T~Ǝj���ϭաyH%�+Է) �����}
u;������/��V$OV�ܫ�	���1W�p�)��D�2I�l,,��٤I7k� (�g�ʬ�!�2���w�:=�\&���VQY�N�ub�FQG'
��Һ��Gzr�RS�|U��4)9�+��g.F�h��5z�wl��5~>����u{�1��&�ybNYE���}:bb���L�jk���'MMM�����KK��}M@	���+})��j�^����1����U��]=���T�dBU	����?�⇒b���|u%��(yt(����x���6��z�Ma���+C���r��)(��=cZ))�Z�a܌���m��uC�)�k�������^AYYYb�0�lj�:��E��u[�����b���Ay�޳���u�wnÌoA@��Щ��'z����NSKK�k�z靪�Z��@t�y������2O�AΌ���,�ro/�c��:�C���R�p�>k�+�֟KKK��ҳje����) ��,��~!n�rH컳��\O��19)b��&���f�,������1~D>2>Kr^i��r/i{k+kڼkvC�k�T=^�k�1��Υ�N$ӯA���Xɼ_��Y�ba��j=sNk�4$�'U4U55��������&���P�F����n77�	�!~� �~�GU0�����{z�M�qS8i� O'�c�Wy��n������ݷw86���'5V����.?�^��#�¯������k�
�-a�������c#���X�d��s8��[d����!���u ���O[�
�7�����a|����<I�|zV��ֻ�!f$��:G<�Hwbvf��9�����?� �dÿuu��cM�A�ؘAm>�Y�i�����nb�qѮ$��H�\�٤6�Q�55U6g\�b�������OO����������x/Ӭ��6���ĠW�8~�x�2\q�=�s����s�X҄m��/�l��\ꉓWR
L:�9}�c�;{|F���7�h�
���1�n��W�n�l
>��S�;`Q`U9����E��6��v3|䴴FcE��Y+C����{�GH�}R��/R
��R�4|A����g�?[�3dԌ������X\���U��=P�n7�9����.;{��칐V000����GGg�(�7�RZ�yט�;��������7r�1��ιX����]������l������ٱ��~�&���!�z����4��q����
[�<���~�b�z��+n#+���8��v�$��ա'ޑ���(�T�A��A��9bU��bb��筺�����[��\�4�$e�s� ��˳¶Xٶ�;uX��0ɴ�v��]O����|R��ìu�G!���x$�z������Z\΍�l�4c�_ǡ����4=�ɜooJ��W-�?[�ݵiƟx|�v�<�^{ 9�������O��w��o�����%1��}�>���k���kJ�knoX��)l�a�2�(K���#�N�f2��;l:�����~��_�0�+�A3j�W�+i�D^��h��r�b$̰S&2��K��'v"9�fE�ٿ=;��4I�j�L��e�H�R���x����.��᮰"��<�ߧ�^��p^���Y�j1:"b��㔓�3�ɺ�_,��}��5TT�i��zVV�ӛ�\S��mO�a}���������B����ݫK�r

��c�Z��V����e��A[���GȊ*��~�LL<RAG������:f��@�T9��-�+l�)�PWǝ/�G<Y(Q�E��C �Mn\417pkp �E �!��/ԕ�V9�I�-tDGF"����	Y~����.�
;�K����{��M�D�(��y��XUD��������(�j(N�nҊ��ve$�"���D�o�8�;��D�T�孭�W��@��mI�`������Q .��������H.;5V�/�t���e����꺌��������������n�=�K5T{��V�}������E,�;m�=:^dP�6v
t�=o�\��+��}F�� ij���wZ
�V�h8�^�~Yv6)�ns�T���/��&+�y2�%$P����F\=u���Zl���)i2+�xh�-��w�i��a�|{���+Qg+�5)�k==�B�^�i�v

h�ڕr4nP��P�\�
6FV��y���Tь��J�F��i��z�Y`�mU���7�
z��a0&

蝁��Gw�C4@��{i��`u�|�
Wg������r�o��U{I߰�~�/�U�s��V�['�8)���Y��dS�#h^%�Z����%�)Z��V�*����;wX�o��( �<Q�*u���Ѭ���;�o�l�vv����W�#�+����ڥ�*�|go$Qr`����e'���N���H4�y��z,�$vHNMm�LKt#c��eg�|z�\S�)���@������.��lzJ��Êxqy:**�؝�,a�C��Z���-���T��1���C��P+�,��£��q��j�гB���������⪜�M6`_�'�v�Ԅ!:���A����+�3��q�-X:�[�ǧ]I�Y��=�@Zw �79��!���۫�l�x8�* ���s���h�&,^�l|=�ջ�#�����3}HߦdN�奭�,�)<^72znSn��żg]~o/u��d  �J�1���I�������[NC�ة�/�i^�QX٤S�wP�g6�5!*v��1X0F�a��<�����@HZm��[.����V*~bƧ4%&�]���4����iV�'�Lw�<@�E����i�Ra���9;��$�v�w�V�S�_�GJ��ګ��Z�<Y�|�F�7!�93�PsL�u[i�o��/̤Bd�2ҌF�z��F�Ύ��{��Ġ�#�Cǡ�n�&���MC,R�l)���2ˑ���8���qj�z~�T���kp9b����AB$P�x��R�$6u��|��R��i�����>���)��oV�֨8�lHj�N����4�2���2����B����V�Ro�6HF)�==>�dll��Ʒ{[�x8ׂ-�d����P�<V��u��]t�BO��������5���q`}���N��z&�~qeeg��/ZQK��FFFFp,y����Aj�GR������9���{����h`�rs��x��� ^��&���ΦT���-(/T�Z� hl�4m,))�#`T�0������ͦ�~� �XDС� ���L?����$�FAAA�ɉ������Mt�h��V���c�o}}o�V"��O�q��瘘XU6�}��*���&бs1�����X�i``�Ob[>���R���x�i�t�>K0�-���ި
��#��bL�7aa��G�eD��>��Vf۽��'\.��-U+�_9�P6��\m���R�O.zf�DP� P#s��Z��5i���,�m(��u��Ƶ�M+��;�:+����� ���n�#�FXR��`v�ѻ��R{o�8������k#,liC��89�Ҕ|�T�ݸܛ��9,���+_nc��'e��TW?�䛹�R ,$�gQ����T�b��j<ssݿڈ��㽳ϖ��FW(t͟ǚD~�Dj�~,[v�{m����ے���?[��ƠdY��rYU2/�#ϪL�3Ì�&�`Ʃ�w�!�깕�ؘo�.ZYC�#���A�ӳU�k��`g2K�Uஉ��kq�����r���bV�0����j���q�Rᷯ�0�LBFxX�<�rZ��=3g�)�/��$ ��YX ��mK	�t#���lV�":H��"KJ ;�ZZFfk&����h�g��92})7���o���|8UC�~{��1N3��[�jI��z���<�%�t�YnkI� H�s�S�(�]zG�!���	�����x��5��L�f̜��B9�4�3�%+�v�x�D`�~5����LAs��oUIRq��y8̲dc�0\��Ɛ�I�o��h� ��,�)/��7��SY)WR	�����hݫ�� ?>��������.d�7�'02��~��̿�O>��bO�6�����Ұn(S���|1h�f�c��������9��Q
"q8��p�ɹXk)P��KdН�:��*��'PHD9���iQ����l��%�Flpx�ǐ.�9��	IH@����}p8���� Q��l���7t���'��_�����V�bR�)1��n�����9��;��F����L<���`/�߅�|�)G����==��~��bQ2��"�1��)�y~p��UD�,��}5;�Q����ڍ����-��ے�4�P
m=G�x��%�����x���Ƿ�x�&ZMAhG�ZJJ�R��`�2R}�e���ښb��\��;��5�{QQQI����o:�ߌ�bj�������)9�C5����͠����;Z��� ��>�&�<K�G̕X�v��0~��� �������[*c�^HpAW��46�Z5Z135���������u�)_]:*��⮜�3;;���y��ަ;7�lwQ"��i��ʬ����O7�5�,��Yt����Ӿ��?<~�\D�vAt����U����1�.q`�,X��/��v5�T�t�P.�I6��Z��h�N}U9�4ٷOb̦��,���ӟ0���q������uS!e���zm�K�7�PF�}�2Rz�Ł��U��:��x�����Ԡ�:r9u��B��^��V\��n쌧qvƐ�W�͘D��b�}��ڿ���=����%X��digV�IX�d�v��ヴ! X�,>xx	ñ鄶�^@��?��������}��_�>Kn���P�PB�S���b��A�j��a�n�q-,�Н0u��Ê�ɱ���}��Įg�F�⢚��Ѧ�+�(�?q�t��'��=�e0D((�$v[��� �e��ǻ?x|�	\�WW��bs���D���b�����x���� ���p�wFy�{(@��- eg=&��%���%�[�����!C�1���sI͋��'@�S�$�WQ��7���}
�p&���8��y]���N���N!�[K1�����|�P�s��`O�NT#i#�;TLi���G��@�4��e��QgS&��j�!���7�������B~��i��J(�U#ft���"=Y(S,��eqAHa�̗�P���;U�a2�e_�Y!�KL�$#����F��`�+Á?5"C�fw�m/�S'��1FG_Q��赛s/S��d���2�1Aʫ�	�?�
�EP3ddR������Ŋ��B���t�rgMa!(em��X�P��L�(�	L�Pl[A�tx��|g~{��Jp=^ŭ����х�l�AE���:��%C�p�q��e�
��%��|��
J�4撄H���F��*�4��?�<±��O����gzv��\	6ϊ�5-�_T�����ef�����.W �H�����V��bab�O��O�ɡ��$q����ѱ�w�_�>9ju��)������������abBmq=�v�=\�+�����n[��ļ���4��;�l��x	��� @���Ȁ�t��g�"�Ҿu�uw�I��,M�PS���:���$�N�������p�͙�`�P�P/��P˅��'����uҷ޾���+�yqRy
|N�hscc�ϨYO� s��Yz#!��M�� �ٿ��Ijk�����)�t��܀�C��d�u��M�%�\� i��͞O08��g@���^���v=p������sFV�9?��XX��;�Ȱss�qѴ�Y� !H���6��lV���6�Q�O7����!�L0M�Sv2��01�4)#��~0f��X���,�2��Fs$oǛ��j��h2w�/�����3t���mC��{��|W��A�~�"��e�ԟ�D�"�kI\�xVf��0���Ԛ>W3����G|RUUMϛ�oWBi{Ӛ�426���3�ȸ�_m����*z�1;8��/p�?�����7R�E��29,Н�VU1q=?��Å�`�C����䶱��	�f�W�`Q���?�:m��)(����Έi�������%�^~(�CO͋��xJF�K��������� x�W��p��H����A';n\s��E��a�$Bʽ����6x�����2|f Cp鵳�mg~�^8A/;�p�WVUMg�3�����E�W�C[*�0���{k�s�ӷ~upP��B�L��׻%��LfZE�?n�a)I�ˇ��/��-��WdǸ�+.�S  �3}g�}��� �ˠ�ڹ<gi6�.#-��N�tR��(dZ��T��: mS'����]8U��-���ƉDđ	jA
x�̸�>9h�#��O��V:@!E���K�%6����?(J�I�4i(B�v%|���R���ǁ�����su�����l�����~w����)�����
����ƻ��\�4�/���,�^�ߍ�/)�à��67�PX�B3:��wZ �bg����ҵ����~�%���D�k-�S��%�֥eeS�c����z�W�f�`�����!�ɮ޽�ڥe"��HG�O�#��%�b�Xo�:9_k���	_6}1�NIK	�; ��z~�hNx6iE9[�wWɓ-��m� �b�5{���I��+>yr��j/�����v!���lPKf�ϗ�r��F�qߙ�'�v^�nq��d\���[2�� +��E�c����V�}�]O��c��;)��+`%��dZ4X�b�����w�M����F�OJ�l���fc���������VH\\�֡Ȭ?�0�"��<@�%�1���`�#��񝿨�	R~�K¸�����!�#ot�U�t�P��P�J�<9C��= ��~�d���p����H��۰���Y��<�%==��������;�x��@�iE��2�S�4�'����w�&hf����&�u�@���J�V��7T���#2֒p�7��bP��X��t���L����˟�8Mv�U���h �}�C��V6�t��m����%�h=���T�|�f
�����z����-��`BT4�޹Q���CL�nB�>B�����6��з�`�﷋�>��ӥT��N��u�DbG'�?���TF�rm���/�@�A���.0���_2�$;�S0`־����m,�M(���Z�n�~�ll��\P�m�TF�N��$?��=(*H�嫪|�[�aN�c�l�����5F����Ia�3�(Ϊ�&���֖�l��ù�p���}��iBm��i�訨��[��I�K[��B���D���A	6�6{�ߜ�c����!;�_Vv���$N��Q�_.r0L�(n^n���=1�{ѥD��P��Eāzv��9%J:��Y\||��\�s�Yr0���D7�Xt:�  X�V��i������X��7��^%�ט������|��k@U�jU�3'G(�ZYE L'��b]6P��z����RHy�?�6x�%i���)��03���x�q�~�����;�"Y���2�("|�ڨw5�������o̒R����CZ2rH���`�u$H��a��⓲÷V�����vp��2�?���4�Rr���E���+��F���7ce�1�*7���L�g1rx6-�L�̸=�Ȩ=Mf�W�s�� �����U�lˊ!�W���Ka�YZ4V��n��#uHy�=�
)��Q����}V��[{�C�!�-�h�h�(�g���6��J��^����[������Gbk7;�K�ث�_P(��E�h��m	���+,H�e<����S�4�$��`N��7��-)�_��**�-0�n/I����X��ÉV�щJ�z�;��)���y������/�ܼ��3�-�����z]x}y�����z��m�$�G�����װ�+�~���b�	��`��?±�333%�qg`hHe�_�T5:��~�ŗ�e.qqqP�k�}1�@4q�3�1�{vhV	�Dv%e��<���JK7���,��D6{�vj�v�auǰ4TVPRʕ[*���>\` |�:�{���cwu�5-b�����amC�xx��TA\�?k��5��ǣL�}�>_;��Ƴ��O�~Z��er����d|��4[�;�_�b�v����NKM��(F�·;'�|������ocUV�, `�{D���u/,�:�=���������D�lll�f�ڲ�mu�eA���|#�����I��IU *$p,�a*#s�		Id���?���Ԅ�F�5M��Jm�����B��F�o�U�4y�q�i��-�M)RJ��iL�h��>2�&��bP����W��I���+C�<�ZUGxGZ�v�(Bqr3+x��-�NL,h��7�H�,��Q���"4$$7R}��f=��3��Hm�WmV܄n%X��3��?(ir�U��MLȫ��q�e'��c���=;WVWg�Fg0QQQ�z=D�p �w!X__����4�o��Iw�g�i윎'( ��[��Hy%���HI�I�
 ��y�S:�t��	``���e�c� �_|?3�Ɔ��ff�A����m����%[*�t㻌���k0#F�"�S�!!�ʞA��;�s%�C�^+.ߝ�enVZd�W;2$�$3�� O%�!�hO+׷#7ϰ���A��7:�p7� ��_���O����P��4*���ibf��zO��|h|�P��6k�{h��#���]��i�rxA{Px�m�[奐�Mppq������}�N�E�� vZ�s�J�m�{�V+�f2V��{��v~\�t��7���������6��>��_��|�����_�t2��i��5���bc�~I�:�MH�xDK���SWE�����B_��O����*lmM���D�='H�9>�D�O�Wdn�<�h���`�!�o1��N��S���������b����o���I�J2�h5��ޡ�8�?^wǘQ�����V���&&�k(��<rB�֠�6�ҳ_`�c�suA���h^^.���� �D��ee�'�����D��#�o<��Z�dD���rs�z���4&��Zq93���1ع��׾|7=���ņ��J�a<`�/ooAkbZY�>q'��c~�AW�j��-���~~����Z'g��(@���5(Q�������J分�^�8��dUX���N�C�
O������E�Ґ�k��$C"����7��Ȼ$�q|I��JFZ`������G�Yud7����ż=�Y�z���3����F:W����^P,��cR��O�!5�"`(^�<b�S��O/�+�P�ʿ��$���Ml��l�5Rt�0�6V�q��G��Pҩ<?����ë�ϸ��7W���A�붔OVn
I#�����Y(�e__]�Q�P2����B��Y.�o���]�94���v"u�=!��v����2F�>�Z�D��ϳ�x@&���`�[��� �����#�[j���_�w��S9wÍkMM,��m��ҫ͢�_Ӏ���2����pku�X�-`N0�w��j-.t���둸�X�\���s޽��;x�} Za�S&p?�x�/O/]��!
�;��AE�;�L&�8��Ulm���#�N��V(� ��ହ����`V6��(����g���|�%8ʛp��B�HVZ��t�Z��En-`;��H��ϥ���z{�ϝ���B�c��}�9`M���C�D(�kjlԛ�ոk0��逸���	��X����q�ݰ�p-C�������OU���ip�x���3�C��[�+>!&��MP`���ծgo�Y���P���������'���I������%�i��@�"E������*�*M�F�xu0�\�P��Å�N@�PRJ���������oT2�l���Z�+��cM	�q������~���s�
QoV����sv�{tOĢ�����O��z^��E�.��mvZz��YD�������5�����Ճ��&� �FN�w������U���&e�! �$�3'�b���G�x�?ӷ2�������Z��
ҝ���4N'�i�Ѧ��'�s%*[�A8�KK$�׮>�~A��Ԙ���+�M�VG���~���$,����_/)�E~7 j���X(��	�FV�D�s놡=3n�B7c�WH���� a�i�t�l�s��]���5%��f
���P`&�đ^=�ϕ,q��˸�2՚M��c�
#�\�Ent�(�rj@�
�	#��i���ONP�I�::1qt 4��_�,��4H�4ם8}���{��ug��b���Hd�F��ch��Ya�씫^�OB������`�JL,;�&�{*�������R����⻦�y:ML����N����yC<�^����Uzk���K������v���C�oA]$����i���\anS�4&�@��9�L�(�����4�H��Fu��4��f&����.�D��.-/���ΐ��N�v��i��v.��?�$K�6X�o E&��^�=+��5����(wڔd�
R̛��Zw���>L�wO��
-A&���0iؿ��k��*��������K����'5����S�<"+qD����P6Z�V�E��i���w=ގ1U�u����D�6Q�X
& T���sЊ��!*��XR�9]�7�c����xo�v�'Me�-��ߡ�)`eE�4����k��hvoRקkb#�#٠
�*"�GJ���־Z{�p���������l��H8����,X�v@�� ��L��vg�_|s���$�(at�2y����<K��i~|\\���!�\��0�|\	���G�Ʃx����Ϗ���|]����K9������y&�y��a�_��%)!���/[�o���}�X5en�!�?��d�.��+}x#A��a������-`��p>��~z2{�=_Ӵ�p���eV�z�����'�4��cϚ��&G�9�ҿ�W�+��&uDX�X*Ŋaoo��}R��L�!&%E2�cmumk�5�O�4RUA�x̚�`�N��,@(�Ll#�}���¨����t��}��q�0��k(J��M����*��(�J��ST$~��z���"#���/���� �:.�_g���]�۳�G�_�#ō�����V��v�37�V[\u���R|I��x�7G� �zy������J`P�(�q�{(�v������ *&"����㌸
������y�9̷j���F'<�g����󥅥e��M�^SSS�j�o�)p��,RB�Z4	����9	������ZY�ى�|o������$�0a;\��~_��*
<<|Н��1hR���e�`��LO��R� �)��2����$�
~�Q�7בpr��ۮIj�Z[G&���̀���m	��n�27��Q�ئh�U���D� �����zT'�d7�����������u�؂��^�^$44����%^xxx��oϥ�?�~p��������tߣVy���t�$BA���7h{�j#a���b����(�ǯ2�)�JR�\m�"c��D6������X���II
5騵���F7��VaJ���Ϡmt�Sя�.b�D�b��^��m�%c��c7�W�T�a���#����	���=و�޹L�VHS�$� ��n�5�~���bO������'U���ǏU�q�~�|^/�$1�0��i$v��9L��P�� ���by�R[X��I(a�P�D}0���b�=�\��ک�-�,Q�S�c��+����YL(�:� �n	�;d��I+�x_�Db����ޖ�5����%�e�&�-�������(A���~���E(R*V�X2r�b� G���f�]_�"Ɛ4�Y�`�i�{� ���Ytfj$>eD���dV��j��?�����8�,�s��@x�&/�K	`/_� ��g�����	m#�l�C\�����i���pNy&��;�u�qddd�O/�脦?3s�ǂM=d^SS��ȅL�@�Q�	��E��;Z���vOz?4!�8nnn��L��-���c����lzЮR�Ե�:P�چ���ׯ_7'�|�5"\���6^�:Hz�S{�խ�@e�#�����i���
����k���$B��?,�������绫�L����L��O�8��*e��x�6�O���5J v���)ԏ������� ��tP�Y��˽�]�r)�A!���;�����6굍�	��:�"	�FV���2���
8�a�oyL*�O�e4/��X�:;�r��X:��� &Á�uN�o�B_Ѷfd�R��y=~#���̫���ݯr����H�y
��K�>o���8�C�����"R��V7F��N%���0����kڡ��*����@��9?f�͖k��^�\h�k���_�\�r�]k􆀾�P=I9��~�KUa�H�đ���6<q�6 ��.��#T��E�K�$�&1���h*��~�Z�j�sJzz�_�h��1�K5v�16FF�.g�Y�鏷5ů'�e�


f5�����o�.Ï-{i�B7ЃnYo�����t"�9���F�a9	��E�m	W���]�P3��^p());�@���8�-�\	j�b����Ҡ��[�ƍ=��eVK���O�'�9jR���̐����nz�qq�Z}��O�:Vˍ���l�o� (((T^x<�iTV?���:6� g**<���y�𽷷wi�v+x�:�,2��oO��_]�_�x���r,�#��ׅ����q��;"E�Ņ�d,)�D��X��!�H
�-`�8�thB�E���^1��w*|H<p<U�H4�о�du#��p2_��dff
��8�M�����[�Bց 9�0	i��S��?���Oj�k7�c���_&�	��ii T�b:.7�ıP�D��Ѣv���u/����x)����233����9�-V���VK �	Ē���4��6YǾ�<+����{�Vy)E��u	��`�SVSU�u��b��⊱�w��"�+�M��|`Y��\���G,b9�,L�������!!0�w�`uF�O���6K��*�^�k����[d�1�߷G��O���H����I���� t�k-��7�99ճ��EDŶ@K���\�ǁ���jLZ���k��<� ����׿�TS@ɠ�& Fͳ5=3cwv�*ޒ[�g�����g�2J7��N�qӳ_�o���s��=nk+��kKKK�ښ���SPP��mv**uӉ��¥'������b��a�����W�=��:=�M��~W1�LM�Ġ��r��b�d�e�)g���l��g���ޫ�å�=����C�[�@�Md@QQQ�sHXD����lO��׷ʳD]5YU99��>�J�;j JY	��OR��dC�?_� ���{������t�ڽ������'.�7!���Û���5�qpG������^*C35]��u��Q�{��4e���S)�U�{8(�܇h����nk��A�q����Ƞ����282b�V����8PArC6�y
� ������t_�'�gfN��p����5�#��%�b
	�Q�9�7�w�@ض����abam��yD,|��G��5Em�����D�����L�Z.��~:�n�;n�ͅ�ut��xKikx��'���%y�S��������΀^���z���h"2u��|��I�i����9�����y��~��(%���=��ޅU��\@F�"��uԛI���e/	`d�.���
,W���cRE�U!�!A}Q<R9|��*}|z�j^�����Z���i�f� �G.=��j�DEECBI�X�_Ԩ�2���H~t���uhBhjr#�KqZO�s��JĚu����<��V��:�ߣ��p��)��^a@`��&f_R9��Ǵ�PPP�n���M!�{� ������bc�e3���M���F�ߧmO�I�越(��iZ.�N숏����ĔH�M�7~�%���vA�`e�9���A��Z���N�A���;��w�Y�:�y4��r C�5u�ir�Z(s�?���Xf�-k/P�H�!`��B����o����F$��6 �«��A�P:�i��^���I��c��^z ��
�:�2dK����=���1�����u��z�T�.lWyw��+a �*M��Fu3*�ML~OV��!�1�p]�.�|]���.�p$ί_�6��f5��oG�H~SW��+�����d*���z�Ua�lS�>�Air\s��J�)[���u�\)��t�����K,�T&���}}}���c�k��acc�o]��^����feQ�6�8j��+\��-�C\[������-�w&P2�++��{�ޯ[Б�s�yɎ,�^B::D&���kh�!M �#���5=0)�m����k�#ז���/��3��W�軃1p�+�m/��Z/`�y�2)
���T��J�6�{��ҿRT��2��T����~Mq4`Mɗ7��E
���GT*�-�N�r-��lZ1����dlⲟ��v�����V��N�N?'s'��gkΫ<��,r��'#�MH��S(�	,�d/�h�X���_mv���*r,HX��%&�v��
��CM_O�~6��8¼�S���2��N�:>�ݕ~<���)$��tJ��⺊�@e%%��h��C�mF̸��W\�55'"�����rv6��@�h	��./d��g�ePqp
�mn��yCoo�F�M�q�p)T-}�&���w�S"#�"�ԸE��04̭���B�p�s�jr����},Kݞ��U���i�+V��JC�:칀��V�қ� "R9�3�KxȠdcS,=���̯CgDDD�(�Y����/��*6D�P_n�x�2��=)5���h���ӈ� x߫O��5?.��l=�L,<�U�K�@d:�C:VYd�b����N4:�r�l�I��+�5��p	��>����v��;m;;F�=�X�����=ӭ#thD"�����%�^��׀��z&5m�kp�(@���������\Yo}�0�þREW����?�L̥E��3dgCz0~����ЂY�O%EHH8g2V�Ֆ�j�x|ȉ��Q�x}��u)�H�����1~vǗ����:�?-f�����IϪ_���
��R��mp���˷f6}�WU�؉�R��{�,�خK69������[�utm�X(� ---� ���tww}��.锔�����3���������s�o��{f�Z뺮=3k4�Ԑ�����L����[�ۖ
/��%K�p���E�r?)�bgՁg�}���a@E��%s|��&:�pjMM��[<8���9O�6K�W:7G�c��CC�n�-��7�G���Y�Y�}�W�Rm3/��Y�6��'�G��1�Ijp�p?�N9��M��3c�=����h]���_�>���l�wMUe��&�D�/�X��X�Q9F=Z��q�ϥ���ñ=Y<�0���'�V��vcR��kh�#��@���Q����N�"&�Р�A�2.)�������k���;������e^��D�AɎ`�QQ��Ml�Jѯ:Ǎ�(Ĝ���O�-<�/�e�B�-������1�k{�S
�]o�q�<M�ԉfM��A�RUPppA0�����#�����F~$qQQQ��t��vn�����q�~��c�Ñ���U4�OG䲦�z�����D�xrr���3�˝1��1Ƥ����L"��z��k�@�h�`�#����y����ovn���ک;*���=e-����௶�MY�q<��^��5>�E���ps���t�� Z�L�����V�ŧ��_1��3	����Ku��#˫��0�q�:�`�_��6G�j�N�*�ግ�3)N�%%J��D`�s.�s��������l&�����tn�L*��(��o�fi���9p��8��+l_��
�P�s��q*��N���@X"��9�b$4�`���&0������E^느�Y���?`b��T��<+�#�7%!SuT0��^�5�R��k�\���j b1���Ƣ�;�9�YWEss3�4�CDX�B~��Qn����P������O3�;I�rL�F$��P[t��Di:T�V�ؠρ�>�FK���S�0�qyMMMd|^%�`���t;]�t��&G���Yb����Z� #���F�M7������m7�h� l�n3j�(cZ���
���m������\����2�B�������ne��ʦ�(ӫ"� �@��ۧ)����+A  %_i����r��ű��e�tߗ�13�@"��Ӄ���>o����wr�M�-66�͖ԦzkqWO� s�C⻼�	�E�t2��p�5�-�Eg�CX���Qt�s�Uz�Ś5v��e�p�4�kpY��fg�p��H1�JMM��d���HZ�~ё� �놬����ET��Q{�'+)*���C�γb��f�dyqy�`)x;Ϋw^���AǜAB?�3BB�ƻ~���s�<0�kt$�{��R9m�{�"��ND%�!�K檱S.,�yޞdշ=&!�������^i�_�z�L���@��/ND/\�X3�G+e�WWW��p8,EB�BQ�V�u�mq��S|�
�o,I���ӭ�Z��i[[[���3��U��h�3����ѵ�=&�Z�
h�􊪨�M;���T��ex)�]��	-
���|*�����M��|�μ�9��(�I��A�c�<c��Q���R[+^
�xdơ�w��S������9T��x��?\T-B%�ë�&|�ؕ0h]܂Ι0""M�GEӪ�Aa;H��4�i7{��1�(i�/o�ed��?�/<�>j�i�ݺ.�z�=��]�����APqtD�=��LIIyc��,����A���w?�Wq�ϣ��'�m�/Jf�{8�~�#'�(X`c!�XV��J�;��Ou�9�Ǿl%��ݦ�?=}8ZBn���V�:p�%~�+���LM* B,���E��(��0g�����fd����B�A}��A]�'�R�aMⰄ����Z�(�nO1E�Γ��,^f�c���ҚL2�!�պ���i�b�^�����&'	(�(A��*�ֳ�p�0 sQAA���pDd8�Y#��[��Zv3���z�d�������XX^���P��������"岃[em����/B���L�B:M���qx�b�R?y9'FI*@W[b�ҜI���+���Q�D�PF�xR���K��qݧa�Q;��C��c9Hi�Ǎ����%zkm�A�`W�T����&�./��G�8��0���
��ٔ�EAo�7�����+֑�&;���붹v^�G��t�1��%	IQ����F��v��sa)0����2y��y��+<��J��u�;H10:��U��&+��1o��R!��־D@@x�Ȩ�ijj�ŖkImcI?몮R"�7�a����Ѓ�L��p�\��D�ϛp���� "�:��.(2`��������ɉHЋv1ܙ���oRT6s�ƃ�s����!�Y��
���7��iX�(���&Q��c��4��h�c�-z���й�>=���X�K��ym���¤� ��160����⫘���X��W��vx�_�[������m���F[�T�,��"�Xb���?cF7" i�i��ϟ�_�:b�f����]s}|R�ώ�:�����?9�D%�̍�YH�kN"�2�-����qs���*,LX�)Z3>��d�����PP��(z_�E`�mS�{�0�c�˛�����>[�\��Ȳ�7��T|��^�����(z�ْ�{�]��Pi��T.�&�3L+�����!!�ii?j�ZZ���{#���澨��7[<n�\�襡�C�+��E�644�K-��]����G��q�����qm��'�WW�˩Ve|�޸t\-&e��w���W��<�m�G�� �h[��)�"��Bn.��l����ss�`!�8�4�{ɠ���T6������I�x��t<e-S���i1���Z�����M���X��,���o�~ʃ�����ӟ�X\�4PHY�٭�P�Q���?����ԅ�<� [n���FZ,������Y�)����1�����&>���lId����c�10�}K��1Z�%	��f���}hc֬A,	�~f=S�a�S6~��9���6���g�
��N��c�%,��Wh��i����x���*D:b��'o���Z��e��Y`_7���Mz� �%ge�T�w%nr��4Ӆ6ѵ� G-����!��YJ�����;?�	�M�<M���9�x�-��c�>�NbU�D��K�n�'+10$;��{]Iu�q�f��m'��*|C��,n��	il|jrR���`0�rm_E�	�_�[�d�h�0�4���쓿��K'�״�����/��>�����c=|�!��o� jܫ̇`϶�	Uk7cc*���t%���^�HO'5h�*��ΥI;WZ�66u-��+b�JU]ܡ�ͻ�ϟMM]���Ͽ��V��H����
�/���n�%��@��D����@����1�q�,���B�%��ZZ)Yr�L�r��_/��{�#E6�H:�ةB$���M�"����o�������|�LR��Lii���sg��\��r���͋��و�@�B������%��,K�J�^�5?Ϭ0ZV���j��+;����BR�fR���<2�?��κ����s��.�Ʋ����?����,�)A%׎GNF������P�������x��=) ��1�J�{\˽[l��whO��-`N���.����L��¢J�E� Px;�������ʺ�٦�ǉ�lN�Ny&�ic��$�f=2��N�����DDħ�\��))�x�->�R9
�n'�}���U,�;�r��Y�W��a)�<=���[[�͖_S�|:���Amg���QZ]���SG�e3+��p�̛�#%��i<�ƿ+�2���Ϙ�1
@�'A�ɀX�|`��xq��WS��Qʦ�lJ�����v]'"��������䒆fX���w�ܭE�6��(��1>�Q�FYZ"���_$��� ���3&x�S���ɞ-Ak�����F�&'���_�b��,�����p�G4��R�3�������88���m��gBB%-�OL�1^�&p��XZ0�ܺ|$?��2�&󵬱���;?���4�[$�:��<ML)&�O,���:M���U����ja;q����^���zx{7O���aq�m9>vH�Z�Vj���3*;��a�n�d�Hmp9(`��xdPc�n�q��\��H�<�Vn{�2J�o@N��U�D�..�4��)<:֖���x�OMMw�=�T�t��.���Z����B�h(�-p�f���s ��KGP�#��|Y/�R�M���n����T�ZWx"�3����<�nЫ��K�m�Ã�)�te����2w�J7/��m1M�+k��'׶��zݞ��|��=&�&P���WT�L���j��}�E������^�]����ϧ��7�V]rŊ�2Trr
�3��o�	�Ӣ#D��V��&lG���L�M�ttPs��3���A���!�h��pۿ��Y��w�[J��v�P:׀�����AS�߿���'D��)(�����X�UT�	^��6yLdX�GFFڹ��jz�\Dn�B���l�
�S���w��XA�ɫ��2��3_�g��2��B	����粎������N.��ch@MmҰǈ>����# �Z:xBT�cm;�j��d������tk���Ub�H����&uL��9���%��b듦sK�B��&?ѓc�%�Hg��q�UcG0󛩱ѿ�F�]�{�����[��yVm�hu`#�y�E�=Xk��h��sl���0�������C�}p�*�Z�L�\E|s���;%77&��ϰ�q$Tt�o��O�ۦ����#Ҝ���}��'��V%�/nO��d����Fٙ�,J������Z�h ��4e_�������z���H0�j2�en犒�9�A��!J�P)���,����B(ge�d���QU����\��jp \�����n����#s��|?�*����x������fo�E��S9��� ����|�4��#c�}��ٱ�b(*��Dg3n��pgB$�W������=�`1×@�0��م��&F�v�����Q���t�ɨ��G�<�\��nΉ'���;�;��H���?v�LXZ�:��ã���>]�&Q�q����pbq�g�F�����bӴ�i�& 0��2x���d�U0l��aP<�ϕ�_K���4���p-�| ���Lwߦ�Z��t��mhX9�z�\��^��3����~lD����APAA��|E,��h��x���k�p�����i6c@6d��a㭌�A�4BY�G4M?�4���^���idV���ݿc���LN�>�w`��E��Çx�Yw�7H,R$�`&	ٜ��P����$ ��|���C#&Ҁ�A�K*Y����0\������%�Y.�r��n���<��ͩ��q����u�ڙG<��D���e6�
iM7$P�0jT�j�8<�Z1
�Q��\)�Y�ױxN�r'[ƻ���D(���P���%B��23����K �é2Vd#�"�۩j���6�M＆�TU_��Ed�S3��$ �u�dY��я;?22��Јۢ�n��mzZg���C��$	j�7L���?d�<�:t+�[6_iy�Os��kx$ k���@��f��2��U$݁� i�e�? m�O���:{�s�ͳṓ�q�2S�;ܥ�
�K�_�^��vI�w>}��������w�W��ַ�a�R���q@���RU>���3B������R.�����][v�y�o�G>|��&H���<,:���R�\��Q���`a���]3����ɶ%���KE�`�k~Σ̰�x&.66��v�gNq�\�P�~Z2Zt�{��?�ɝL�y C��� 7���RR����B�z1��]���Ў��tN�덉�
ӏ �:�Y���i���=���0xv�^50��I,"����U]q1�|�5<�t�'������y.�ۉ�y/����<�%oT�益r���z��AF�A�J�b����;ո�,�M�~9Q�m�u���>g7
�#���;!�B��Q���{t�G[K��浪�ü��\�D�'G�B��9�k����T�!�����P����u�����g���l�ͣ�H��z�:L�σ�,����Y�2`��s.���C=�:����B�뭮�A!&���ѡ!�H���V[>�����g�߁ܖv���8g���.)������d�Ŝƶ��vMj���χ��~�T���nEw��TGx[�T��+;�4����-��{j}@��R�F��{lw����W��yĔ��e��;#)^��U��焐�7���5!NT�l�!�F���ϓ��֖���(�23�E�`p��Dz%A��4��6##�rl�q/��LrZ�wbQg,��f����D���d���lJ�a����+��|֭(Z�vyHv||<
?;55�X����������	D��_��[�e{Y#�� Z�����I����n� F}�526����
B#-�I^�qoBKW�Q���@8p�u�z>�	D)�nr��'� y�����ڴmpJ�%�@����F�QO�Z&v�o�f�ҍa�-�%=���|{��mra`t�M,�����3j��Ń�,���-���������i^������e55����V@���ӳ��fZ2�$O:Q�-"/?h�CDL,s��a=����&!-�=��ʏ�"�B������y�%�c�{G��b�m���뇩����*m�F�����^�444Y��&��F���_�����G8�op�'��4��v>�i��d:� ���xANX�(��Ó ���\����F�E@�Θ����َ�3���{�_ �:�EPK��}}}m'�wx�8��}������9�9�8*��_ck�oxzy�T����SU�z�B��Sn��OGOߞ:���`����$���������nw�jEu����;R�������iQ��>>��Gۗ����wװl�"A��b��;������ ���l9݅�g��*{)nӣb�K�{5�3�/����>r-Pg���С����n�=mt�K:���;����H����<me�Aee�Wfrf�EE)��`Vb:��l1��̲�����ռ�Q� *nk�x����2�A*K�iUAUeA�0<����Q(��T�4�JB�sZ�i0�~��54ɦW(?��Lм�hXx�(k���E�v؀PM���������fBg�jG%lh��k?�����zTZa56sm�8�o�B��t\���ߤl��S��tm�a�l�<�f�+�Z���p6W �� ��@�ժ|��@�3+��h�e����.�����xB�>����d�������o{ٓ�|.��rB#����kk��b��+r�<���v�Vn��6s�2�\�jBwFwlE���ۙ����3
,hi�_�V�����<@��Yz�3w�h$6���q2�X�L�,1#v�sNN���d��Q�{�Ue>��"���2�33���ʈ�fw�} �t�@�>b���n��Ny,����1���Ӫ�Y�A��wCp71�.�U�x6�� �k�h7�u��1��㵼����%:�3�]��]jzz�"����Yݍh�'�K�蔻l@I����PI������FU����j$�����=͕=�+C8t��;5�0��V9����̣�Aឹ�c_'H���>j��l]dSF��T�X����Ӳ�L���k~�u�2V�H�3���~�J�������w�����v~�scRgw��\;u���4-Y��u��67���lW G�po�����r�)�Cg\����C/ʽO]��,�H�T�L�ڵ������f���ӭ�K�[���(4�nP��ȴ_j�X�l�E�,/np�|@�O�B��Y �b�FT���T�b�������be��SD �t~e������n�J1GMS�W�����&ˡsf�l�/�k�ߜ��no�	~s�7�F��d�B��Ω6����;��4�g4���`�ﵵ 2b��j���+v��P~%z:�6qR�GZ7���ɛͤc9a��O����Ԛیn(�E��8�ߴ�����5ɴTT��w�b�&�3�xI:����tC�g��D�������`�2N��-�l���3`�ax��SةUis��ct���;A���O.n�/,��\������ޗ��#p���o� Drv0�}AV��7y,�U�DXᓧYc36�fk�{�Ϭ�_����E�)�a)��*�;�� wÀ�K�g7�����2�N�DܗJt�=k�u��-n��|�Y��,��2r����7_�N�I���:QSWZ&�����ҙZ�vvh铥J)�$��َ�]�Z�g]��oUs5PU�=���������^jQ���� �s�{�����>ɛsuʭ3��j���w��Wf�S�=�a�Ճ&k���,�
�#���Ւr-&�T�Ծs�U��O/�މ�E0�+Әy\t4եD����X��{��|�� ��aq.e��J���k��=���߫�["�7��d%�?z�F�;<�$*���P����g������=�0�t��I��[&�b^FF�\,�|%��?@�Ѕl�ߛ:jWYTuL����|x?s �]/��솳���&(�za��ug�1����TI��MڦV7��^mVT�it��V��wq!d��/l�pd�j蛍GV�2.Qk�ʳ��u����g�N�;`�4���`>7�v�p\"�ps|�촭��#g�p����F��$�!����ZjXC�\�l�/�m˵��gnRx�u-�`|$���P������4>�P���B���4��gʗYPVP�����G�S�4�Y�q�r���qp�;+�&�,�cڤ��ʬ�Xo��dg���*�jWgy��8�g?�G�S/�_��a�-H%RP�%� �D>_�ϟ��W�
��G�+;^��F쀃�6?<J�,r��t\����OE�czyj�h�u˭����@�R#S�|N!�K�<�� �z�5C�,Ǔ��ʼ����H^��f��y�omm�fbw#�vO����8�(D7��=3�\����d�6A_~��w��-+�0�ig�Q�9�����2�4t(�Z�����>"~��;���Q� 943J崍3j:%IRrP�������I�|���T%��f�C|%�6.6��~
n�o��A.�O6(XȄK-�QI�?�)�8w�Dj��}�cA� ;Y��M� Ȭ��Q��x�E��Ф��{j*���c��mӔ�	`��a�vz-�;TPe����$�v�-|\sҡ��XzZ�䛋���8S%`l0@�QB�o4�����\��w������	��t=.(1Lڏ@C���`��ܜv} 5��q�Z/�kRRn{�P�\��q�ӗP�ݗq����||�/�b�-�Nē�[�F���z�4jɭ��{�	��pс��xI�x�ip�*���M��<]999���Z�'�?K�ཾaǛY�<��[dŠ�7��ÃO���l3�qx�do�Ս1�
ЉSaP͉פ5��w��
����*��766(��=g������Y-Z���=��Kx��������pDN߫_���t �1�����H��e/e��8��b/��H��	�a ��lh����0|�s�:6zJs�Y�����n��E>��fa��E��2������o��Yd���¿`g�3e⋩^�� �x�Q�uw����Nd�� ��m1,��47_X��J�9�
�p���aJ�&&i�0����E����n"���v�	�[��i�Ƴ�dh9F��5�7)�y-?��缽7���H���<.���g��A�w3?V�&^-uJ6]�(�nU�75)h ����$v���T.ޱw�ګ��2�vo�ʇT^���98x�����s����ٶ�p����!�Ys��G%
�Q��a��{�´ܹO#���ٳg��0�����F:#xa������.��N��kj:��Δ5�.��FLz"����F�����"�
W��//����v���GF����܉w��D�}���Q��'��ٯ�B0�60�K�J$��@�B����II�Iu
>>>Ѯ�@2���ֲ`#>��ۓ�y�����n]3s'��`�FWb~�?+���2�����ts�A��ž�F��YR�x_J��!&f(<
���|�f`�״���1~�d2�����sч����S�\���Y贆"���Y3]�{x�U���¼�Z�s��dH��?^��ǆ~-I �Yi��%��ՅW�Vw�}b���{vnc����;��=m݃�\�_9TT���:s>���E�p���$��z��6��
��f��Ғ/4G�M��l{��<��4����Ӄ(\F�_ccc�/If[�'���J�v��⻍6I�&���\\�x��@�k=�X�K���^c�dq�y�9�鈒�'ۖ+�o6O)K �O�G��TIңb��..��G7�#p�=�� z��m�X�q���11������ޞ��o���q1���bF|�ҁPψ�##���sX�榫x]�B�i/I��Ҩ��_�2���_��l�/�����.�g�� J�xu�x��N��
�W3�#��V(p������N7b�㦛S1���C;��|ެN�`��<�K��~s�����oq���k�����%��� A��*���&�-l��ٙ�7��;U1Y���]u�I���q���>���), 	��f�73ZQ�L�B���M]8���8��j6*�'�n�����S�_}}}F-��T�7곝����stC�kN�bNN췄ׄw�yEE�Sg�����f�wR\w�;�D�D,.�qs���Ohk{�M���Ⲡn�F�O��tX��鵕���FZrr�2���WMq1c&��|G�˫�wKF��?�4N�u�(0�π����pޛn���\P�j�uX��j��w"i��$�[j���E��P�nu��#.ݧs�=��fg{;M�zp���:܆�j�ۢN���]�V�JqaZ��X. ;�SM�gj�H䀬�y�Ze���U�/�z��6`xSm�����+G��I�����7_~VRRz�G��3Q�K'Ä���Y��.�"�0�=�OsB(3�>���RZu��-w*�d�g�a��Ae��KkkƧM� /iչ?�9��|Z'N�{N̛pz��=ٟRl1CW[��Zy�3�ƨ�����c-�>t�{2�5���:"ݒ���[1�QЂh���M�:���	����@��ٓ��?1��ܸ\;[-�L��������,�M'ה��P�p�x�б���u�F���o��J��
�v9'���H�e��D�z�>#��ϡD��������Ww7�,����o��7�����[��8��#���RPR��Kn��`�]G�w�^��E�ӣ�ļЮ�d����+���]��>% m%n���KЄtG�)��E'=l������|���⑲׃��a1�R��8Ov|���'��D�nK˴�̝t�� ISZ���� #'�v��oii�Б���2P�����|����oy���n�6�����zz���dy-?>��E_���gCB��;k[��"���P��}�ޛ�4���B\\<� �L�&Fz3�3�L/�c��IH"Q1��_�|����dH�D'f/�tqطU�݇;�0�阤�<�̬,L�Ǥ���||;Nh��L�W'xeG�����uX:�k8Cw�i�͓�g�Ֆ4�LOҽ�C:f���WDo���l[�4�e���Ǽ�'��vV���;�7V�v�f�p5����F�2 4�I�Z�� ��$s�rpr���c:�|�u8 'JW)���a�_/�g#�����+������_� ������7��&���G���W77+�����4��_�\ѫmg�a/U����ÿ�"w0з���.vF*T566����Q�8tU6]�ߖ��B�7^�±,S9�Դ��P�巗Tŝ�H{��35����?�]b���Շ�nnu��Պ��fV�6�cx��/�'����vww�陳>f�)��56�3<8��䐍�aQe6����{w�;&���8p�k��K�w""٨����k�kk�ġc�''� 㵵��l�Sex���u��/�����Q}���""݇�Z���4F���7$6%%P�f�;+�Jy��K�us�CKg5YFb*�L�#�2�h��.x��J'�g�2=?����E*�e�/9���X�)���5�a�o/Ө��v]���4W���n���s=\��mθ+�2NZ�{�-B7�&"���'s瀾RQ娕{��,43���4��|���{��y�L4�O�F����^�O
�s'�00��p߸���64���<>�-Rk&�������7�J&$���S>���F٦�'��J�����}q�2�A���"�t�Y�m��\�G�����ˬ�/�̒�������0j�$�)�������߂]��!`�DDD�~?Rz�P��$W����6��t�E��t6�ߥ�Vdt����fTTT�շ��t��>R43B���6�����)�](��H�p���d�}'K���R�����A�J;��^?����nmy0ᛷ�ɐ �;tu�����6&OOO����"]���]�X���^��	��x%����u�������-���hTQ��Z�-L���omlJ@/S置��-�?]��J��p�_��밖T�s@��� y��� -ߛ��
���2ig$1�a�����qx�X�I��s4�n.(��˦�R�N�wM��M���j�ccê6���b�[Wg'H���EE�1pqݎN�4��3������h455��Nd�GZZ�7z<����	mx���o]R� �7,��r�������R�1�F��A����|��v [g8*a���뭴�]fwD��+�:3C8g`�%-�ׯ�%���ϚC8�*z��[
#V|���9��99G<r2�IH�d���^XHo`�@�vBd�`�o��֖��o�55@������/������w�vE~ �q4�9������F<ݜz�e3+��\�F��ð�<��۷pmmm_��@U3���eeeX��@�(�WT�8I���"F�E>1+
2����dh/��y�:ƙ�q	������_��u� ]�s4���_�<Za>���x� +���?VFCC���J�'K&$���珖;��p��=Ǩ/�Ffs���ʕ�ETO@�[����jJ
�0$��͐�]@��`�*� Żn+M:�WtA�-��@�z}�}�o�� �����O6�sv7��F��0C?�p�u��Q@��حF_X�TuD����Cc��5�tU⏨�dEGL�Љ��)��&�P���&V�~wĶ�y� (��wy�i����w��..��_���n����/ P��sP�Q�6�6��,
_�=;6^���������MIIAaJ}�Ow��X�3�ޔ�}���>L��,���}�=��W$@�B7���
��i���D��f���5�P����s�����d�w�	8,�\���	���a�!ƻ3��'�c�l�����\
�'U\aLR���z�.�pr�rD �!�a�|�;s�������w��x�|�^ a���dy�⧡8�aa�/���yള�w�����-���%:U�л�&ɕkg���DcE��)�D���ax߅�P�"����ii4~45|�M�k8G�#���-:FPcW�a��<�.������Zy'З��ܯ((���k+�'pO6�
	����hňƐ�������� P����񏈐d���+Mgnk�^���!I4��'�W�5�Ш������/5��:�X[Z�u+&�f�mp�΋:��iLd��v�3d��gO��*�~���u�H�6<�Y���=t�n��J0�mxaXX�t�৏����G����\����4�q�xW~�Y���Jһ�n���w�<Y��3�۷z�?���������t���r�����ƅ�.Vn�$�f�|I�vy��9�͖�x_2���ݛ�;�z������oH|Hْ��V��ٽ�����{O���X�E��ԙ�#����O��/�G�y�Y���CCJe��	����%�����K$���ߚ`6X�n��0КBI
���A�l�9m=��I��xL|Oԛ輫�j��ho�
��2
P�s���*6�w��3��s�P��6�=�PG��h��7���EI�6���c��b���˿�q[@�F�>t�6�Ŀq�}I����g)5+�K��P�m U��
t�իW U-�}||DE��,,R	p���݀�M��6���J�1k��d�
�zxdiJ#�ʚ,��5(�DFF��^��,�BOK�z�kh+�з�P����ї%%%�{�����^���N=��#�Q$~~~���(I4�Lj��%�V��e��t� �u[�12�(nM����I����K�h�����7���p8���#.���\��d��mo������Y!Ao" ��Ѷ�������@��
,�7xy����NVV����`�9����w,F)�}IOg�q�B8im#7�<"�By�ZSP���(�Mo�V�q�<���`�������WQ{r=����KrCyy�T�j�d�8�б8iS�H�����*��C��"��u]ZVRX����hS:��c�R�5vpdH����F?q~�2�<,� h�O޼@��������;/ⶄ�>H��_>b��X*be?r3�,E�����۱w��G,��A�*��`���ֱ�����1�yiu�3t4��XDA@ZZZ�n-���>�4@,2�Vn��N��@�
�֩)u�"�G��"���01i�S¸M� )7\�v: �Dނ�!�#����L���U��psrr������Y�������u����ڪu9H]J��G?��Z ��/�sb��s1݃�];��u�J'�V��?�����I��͍���a��� ڟ>e�g�s��>kO�m�
���%���
	x����M�itt4��gO���i�iaoL'6K �
X"����M��[S��+V*�@􈈊RF��|��������~�.ȓM]��!�Pa�Y� )��dy6Sv�Ԣ9�5��K�@S���ݽ�kG���8��WH����pn���:!a�	^��z_2�
� �%�~R0�������ީ��s��8[C�rd�sձ�oӚU���1yo���Ɣ��^����,ɹ2�����\6 b�Jm���V�F���4�ROٖ��~�=�ӊ�w� ���Y-%���|�H�P�c�b���[oF�ީR]�Ƴ��k��UF+�¼Z�1{u2X�eZ�Q&����i���%	|�L��
� |fU�?a�`i��h"""��|����*��( � ��?ň���,i���?xKAA�����!8#n�q6d=�W�4���@!�m�4��G	!��q��o�F/Y�^S7sFX��ζR�9���s@��*ыg�8�A�����v9�*�l�#�NgI�P����V��$����92�0AB&�0��wVjZM�9*��N �N�@聡ea���'Ŷ���'po$;%o���+)ʔ3����4�wu���_��Xͅ��2���~!����M�AB�	�����s�tC��p���Pf��;����*y{�Ma���붾�<_�ZpGJ��a�vg����k)�dA��Tv�J�ѧ'7h�@��UWOħ��m%#�*�@j�^Fǆ	�A��<K�gڪ���)X�5�WlTTTj�N�_�H8��%��g/�!���ܲ��[���c�N4�m��2F���� �L̏j�b�i_��s\� �������%��j^!�c��,W�	7==}�ms�^��Ix�;
��L���oJ^M�D�~Pƚ���026�o�u-Lv�d��t^�}⍈�����&�އ�zF�4�=Ж����.P���I���+������	�f��0<�w�¾�(�Z ��Md{.����C����]jo�%�t:��
��Tf�jq'���e�U����S��E����v�d���oo]�J��ɡ�@�DK4c��ړSS��ߺ7�O�� �*E?`{s��A�N����e�w�F�1 ��&����dάnl�p�R���f�x]JB�6ۣ=���'����1밦�A��R�P�I�t�mTM^Sք�[�Y�.���w�OZ'��T�2�-@Eˁ��v�.?�����2
ٲ�A�^�b�u�����,����c@���j��*��D�!{8T��'�矆��\��	�jj��֏s>����������:ա	�
	�"��-� ���9����t3��`�̻	�
3䓩\x�i5j��ف�/�]蓁a
��oC�����(;މ]G�/�G��Ti�_�4��~�룽��n;��is2�����}MH�J�L�ii;�*L_~���K�Cf񇺺:� UYF�P���GH�.F��{n��PW	��
�]x��O�P�a3�����m��s66L�����KK�cא��n�hZ�jpa�!�U**򪱑�7U OE��h�����P���Ђ��W��� l�Dw�{����u��;łw����0���x��@�����W#h��7�V�j���>.�Z0�����Y��p��)ާ_�^S��>Χ�ʳЗ�� �C|-��m����O��R��ѣGf��Y���?~�3�6����Q�d3�� �w�U���.��6��ӪwB�ac,Wzd�.S!��X�h���FE����������$s�@�SVQ	������Dz�ڈOJ9 /�&2/g,T��Z�Ɗ? ���_�N+U�Q�X�RR���Dd���I>-�&���)�>�Ȁ��ū[�rZ�#���z�?U���8�����n"��|�FGVd��y� ��#�G Jp��*�#��TJ}٠�����ؤ�7�w�iݶ�D����?ʲ�C�����~�杪����zb؊�9���T^7L���t��^�AX^��a��ByF/X���Mɠ�E���gl\\rZsR?\��$%����-"~�5;;��ٻ��iM�o�s��&LKAZ���O�6,��9�			���.�i�ZH~�/�f��'���ݼMj������uNNx ����˗�k#��.�Z�&�J��8��t*ԕ��c��:s#-;~���h	���󉅮׻�����D�M����D7#����ڷ��g;WlP �x���O��"� O ��iM��C�UT�u]��n)����i��n��.)�ni���o.����{g朳c������X!�s��R�U#}uyMb��$��4�~6��60���NoK�������-@�|��D��{ "R%�E�{��d9QQH��#R��v��+ggN�-n;cd�Q�^}f߀�v n���Vy���bҳ;0{�|�|���a�3p�����
�d����4_QF9����»��T���E����U!(qd������2殞��u��s�<�	��p���X�_~��(��F�_ݡF�O�X!�Qp��y� _)���\lV�F~~ua�\����#.)IJd@�D�ʝ7�c�)�&���䄲,1)�m�������)8��kF����oBRRq�xvFz&&p����Nȩ�`0׏..��*���D��I�ґA3��z#gp�!!�M��X��u��B�	f�C�6!͜��~/
�R�;.��4��2ƕ�U���F�*�-�^��ʶ0@��nQ��Ɯ���z� ׷��$rqu��(T�b�<�)+c�akc���L�5+=U�0�l	�k�;bu��Y�ϱ�^�������X��j��'�p¤�������~:ff&�;͒K�����JHP&����;�9o�$ڮv�9]Ūy4���#ox1�.����0oW,c� !���?�$
���\{��򂙏/���b9d��qi`�5�ê>�H��̽����W��{h�577�B��/�
(��h�,�\��т���X�<ɏ��@/T?d�Y3 гx���������۫�J~��q��S���ny-%��@Z-�������?*^��D�&
�l��-P'y�uj�����#s{����_�G%�m�QN�|���pλD�f$i�n0�ޗ���M�"�~��ٷ�"�|2%�1FD���:�������ϝkjj���МFC''�NQQN��MaϏDv�9�T������9�ɴ�����z|�G�d8�R�g�ws��j����r�a�@�(��o}=w�'ӟ,FN8��� Ϧ�ch���m�'��:� ܱ���_NC#$g�lD�:Sƹ�US��bl'��e�=�� 9ʜƼ�f�oh�b��ԲLv��ggf~��^U���� S��;scm'�@͊	�sė3n"���5�0Q�K^��àK���	�����<n����KG$�/.�B�:d�����񱵢�1�@�K�u|X/LؔK5����^薓�ej��[�&'�;���y���L��MFX]-Ck��jqss9l��oo��x����4�o��6�w���a��f������ׯ�Q��5����&Q
�@�*��M�����Ghf�:j�gf�c�������. �A+ԏk��l���~�x]��3����� ��jK�pϓ `g�i��/����a;'�?�C�6.12W�=uZ��l�$%=��`d.!aW��ȄuXZ��9B(���z܅��㓓��+�#�0#M�h�,	ډ<\���g�+�C��ބ�"�v*��d}lMI�@!=S!&�ȁq���_�0��s���ܩj�R�d(�-��S�zLQP��"�q�#���g���p�dvC�Bb��
�+߾bڐ�h�C�e�塽2LN5=}}��+h�?4�>��c�����ɮxr�S�YuԐE�n���ͻ)I"4"���q�'$����cBBgё��g������y��EL2�������������Xܹ`PwFO���}1?��SG`?�J\Z�����?b�ڄ��CJD�<)� ��T�{MAp�TXH�����d����h�M�y`1})�ִ�����yyB��Q1ř�����>ӆ@�����*�QE��j����زΥ%�M䃃��Ώ I�����N���m�����>"$���)��8��x���i�..F �|����L�wO�/mս��Ɔ�V2ו��������A>���Ŧp�[w�v�#���x{_��{3���kt���h�����C�$��U�/}!s��v4=�v�x:a��T��/R~�ڧsmcCWV�o��<*
5s��H��	))"��x""_�kQD�DA*��Ύ��wR�LJj�7Ue���������'g���iU��4��r���Ծzlz���f�5%�n�qK��r�f$����G��֬�
�ٮQ�dK�����Н�y�|k􊌾#�M����!c��n�p�Ma�e%mC /���~��#cm��đ��F�����Gs���hwcccY�)J�RL��I�Ur�Q^����!c�Ɣ�onB۫Q���S��>�r�������_�I�L�O{*1L�Q@ �3���\߷�6�݉L�����ܓA_c���1�*����Vi���<��e��� Ĉ��P�fy�6���
s���a�N��L�dL($�C��?�D:jt���UIq[��~�p\/W"�L>�pکә*������i��H��k��)�`�54��cb���^��̀�EKG׾ ����ly���)�߸ �m#/﫠������L�h�ʳՖ�l�<��H�G?ɱ>	|\I	���k�2H� pK�u*<��h.S�dhXX�b��r�=��C�����"�(P&�pr�(b "���27��UlGI;Y_X̘+c�c2��j��:����h��x��}�o{u�������׿��lmm	HJ��0'J�̼J�47�M��������>;�|���������py��RHP�/x>mh6r� �#;�`���0�t_#�h,1���{�:�����Ȝ#d��6�'C��A�|	\�%T��cGXz)nZ�V�����ZaV��;��RQQ�l(�*�w�P�8�V/�''���w�ˉZ��#���iQ��7�_�i�! ����`�9�ٱݰ���_�%ˮɺ/�ǈBJ)��Rjy�S#�h�h넱��XT
 �����om�+��m!��	M$��e���S頌R u�l,,,N���-|����S^&&�"$��3x��q�r��M���3�x/,hC��x)��R���$������2���)	��+g��k���Y2��kiYc01k�Ad�r&1&*��L�}Z�J�A�?icii�����0{ޟb�y��r���� �O�13��q P�?]A��"豲�BY����\T�^����N�}t�$j�b�@v�t ��R+�g�u5�����6���i-�m����Ţ1'�>Ev^+ϛK=�
q��R.o`X�F ��&��U� ����|�5j8>��FR�o�U�Y�����Su�,�(�j��&6�, ]�H�}{9�Ο����}=�U�ՙb3&.���㪍��$��%��ǑqqP����쬵��Fnn������������R�L�3���III�c%�1�J�+�&AM�C��Z��t(0��7����cOܐ�f������gb8pĨܷIBB�1��ޥ�
�gr�rvJ��
ƾ�^\�=1�:�_����������j���huӊ$���
��+ͱ�uq))_�{��)��\خ�N��ZpĲ�bW���N���R��biTZ�^ו44����`b7�0���7�w؛|�q���z�x��_��]���8��<6��ԓ��p�_�B��h}�W�=��"��!�[�44�%�����H�mlЂ��?�݁�FE%�h5�����}�S��ڈ��"]�s��y��������/_M-%��U�n��H��un�����=��������
r�"���'z���ふ���ɡ�0uDD~c�q%�Q3o?�Q� E�73�4s�����n�a��P���;`�cm��0f4��}�%A��!���������7�L��M��3u�H�NJ�W&�~z� I�J#���UU�r�^��E=ym���'�;�:���o��000��̧�v~h�8�w=�[�h�ɚ�N�PJ��r��`c����ƺ�2W>���޳y��v0��x��dye�w��HS�H �D�6uL��0IH��s|���;_�jA�_�����@��aaHs�w��X�An��t�ZP%ʻ_�1��+FbT�&J4����==�w��ţs��ݜ\]I��浶n~�rww�IO#*$�r�muuuJ��B6�ni���es�z0T�X�E9�D��.���� _	{��0����.���xyC?��GFF�zL$��Z$����2+*��	����mmmM�1�f����$:����צm�O��dCuV,F&&Ԋ�&���
ڣ�㐢޽!�Z��Á;;�"�:�#Ͽ�qpp������Cr�������]4��pc��IQp��'}�����æ�TM��&q(i�2JJ��y<~�B�@���)�<��{�ɾ_���g,�����:�W���ީ�2�Z��g�0�r�)U���+�]Il��<��_���m�$C�o��g��o	I�?��_J�����KC�TQU3� ;.�fe�Gg0搢	
���5����EY!��ۦY��o������eė���P�����e���J�<�~W��	�o�f��^DLc���2�|�aas
��#{�q�*ޛ���U��T��K�6< "������✞}k��j�ڝ���
�R�? ������I��b���K�6)
L�5���N�,�������
�h ���, p��V$8&�Vj�����U��el�ٺ�h^:¬�v�_V��t}{���fS��5���Jlq��B"���0,��-Dl��c���D������*��/om���sj����#%���9���Rl*kjV��Ls�J5Z!�_�g��~���;���0�g���Xe��������UC���v���a���(�(_�A���Gϲ���[���E%$����5
y����/5ؐz��[��+Kt��bbkgG� Mo߂n0m&��o���Ȋ������h㊙��YD���|���l'��W}�4���k-���բ������R�ɕ��(�\+Y$)���`� �)=����� ��_�ZTX�ԢN���׼%�-�fot�J���~���c
*jNK�Ko0\\\��d ��ӝ`ǕW�֕�<=��D�Ȯ��<�%�Eld� ���i}0_9��q�v�H.�9^O-R$ 쬸耒�0��8�������%��
c�2;�S ������&�_GI�?�C��șE�����iF7A� �$k����hi�2�Q.UEH�O�jjl�,��E��:��==7�n�[�.�� ��[dn/e�[^�����*���6T��9��e0\T����MMW��G�B����M͈���&B�(6u���4�[ut�*@*�R!IT��9�kR{�!��"	:�^��ʴ�?}/u�M~3���*�8�pNJII-U��X�F˾������h�[^^V5!��#����y�ਦ@ ��5�x������k���<���kux͟=G��<�| ��`�?�{�ܖ��a�EΏ����&���륦R?����4��`�5�%a�S�n(�J�t�.xܘЬ�$<�@�;G����Kw�����r+������Ƹve�M�M ~A[i4Xߑ��L�$��Y���2h��B�ʽ��?�p������<��^ #���#=_�z$�W2��$<���t��@X�0�kW����_x�F�@׾�`�R **��"}æ��%�):���j�����ȳ�/���)e�އ��W,���V'b��,�(ѣ���������%�&Y�D�i����UH� L��P0(f;�wi"�����\�67?����9t~���Q���M���ʀѸ�\�T���<��c������[��A-,,��t�Lu��������y�+���W4��c��C+��t���'��?n"q����j�4$�����������ABDLLA��|�cvmA�&h ���˨J�Uo )ao�,4׺n��P&��d�������l���L'��K ���I��23[�=' ��Q`C��j�4 �0�wǰ���a�r*1�'�A�B}+�A4HH�k�(�c�o��6����72d���������F���$��i���H�t.}u	�4$�}��н�bv�\���q�.v�zBHo�,#��#�rff4��ﯠ-衞�x4xoF���')��4�Ã��_�8��mw0��h
�9 	�*�/�s.�,(��utgX]ճ4 �&��e�����Ucm9"[v��H��h���5�%ț��م�d�����0�{��%C�Q{��½����N�5J�(s��d#+�V)��)�jjr�bb��C���裶��,���b�?Phǒ��gms��Y{��t@�J�P����!O�fHR2���`�ʆ��s�=�KppTL�*FV;�J��Q�w�/_ ��;��1'�j��j���� #!�]�g67�ư:��t~g���D^�WI�%F<'' ��^��Q2 D �iǤ0+�S7p�p������G��3d(}����?m	�/�_��V����?����È��b��C6&&ow�:|W���!��wb�I �ł
y���5i9�u��M�\�B֨�fz�]]]rZJ��f������ �Y6cɯ���%���+����ʒh�������Qxb��W~�z~^���7��2�u6��ػ��mmm�icx��u�l��Y9����	/i����w<��(�v9��(�@j��Ba�&���.���̹K~"W<d��%9	U#?��Lo䵔�/��߁~
g|\	TA��Y*�<u��Asrq�(,���f��y葈1����� zϪ��Cd�Mwj��SUU%.)����)��5<::�q�X�R��~A$���]ny��v|���������E	;W'�x=33��Y�]��.M~---���q��Z����.i��C<?mȚ��/�ɝ�<��r�����~K� �שK[�� �}_Щ��Vi��~(��" pZce�S�>>�!8�`�0�ng�~fjk342�V��2��w��tDd���TH��?��gQI@O�{�0Nb*.X�xo'd�)z��)q�C)��W�pKIf���_&ğ6�,'W��N}�ÓTT���ʙ69h�P
�H�8t%�Ba�5�t;�~�$��@L��sڡK�Q�h���-�5lb�p�~w2[@^@�l�a-8$X���ܣ��� �{�t|U�(w��(w	Ro���o�[  �С����j��ޟ�����	�$D��eZ�eSC���{���< 4���7ŀ }*[�x)�b1Y����a��Db.���*?��r
�RMo� ;�GN�ӓ���4� ��j���i��
�޸�����>@���;�B��m�OyDpL|�3ź�����*^Ը�8�8���C�ɖϷ���}�������M��c.6��G����"F�? k(���KLGv��տ��y��g���ӷ~��,?'�D��?e��V��#C胷 \+z�墘��<��W� K�9a��k�?b�0]Y]-w:������I�ٱRS�Ť�{�f(�e
j��� ���5Q
P�	����J�`^X���1=W`%�@"6�����h�g�?0P<���3��A]�^��7ͬ�+���X ��� 5: :	�cB��*Ő���=a`>;"ώ �W��~?�B���֏"�����5`���]�"{8K���Ck~����Jn��X� �}�m[� H8H�S�2b<# q����|��Ą�]wg���tE(b}�tYDh�_ٞ��`�w�UC���6�ș��>Q�Y�to�4�l�zPe�V��Y�v�r��������Z��z
(���T��\��>�mJ�<���+k���BH�����Q��f�À|���i�DX���s��#BM�aEBC�.����@.������B�f �&1���}�8;�h��O���,k�j�Pk�Rィ���g�f�|?7���-C��u�/ʲĴ��aR�� ����9���^�� �4t`sB�LPޚ����hzLg��ۑo�"����'~��N��N-�<I��f.Ƀ\` �f�7���h�_ *�� G����ъm�����I�Gpla�H�W��B�H�Jt�؋R/7L׿�NC?��>��"��4���Ш���C27�abL�)�_H�J������yJ�ŅȮ�##m=7b
6h�Ԙ"$�œ@�p�:��F������g���,�?}j-�5Zlr&&T	�*��?m��5}C�d���ՏT���@���ޥ����b�nD2Z��ܜR�rhq�p)����Q�4�<�0RY���c�)C�����1�[��$+R�� �fgo�e�5�W"blL�Ζ��-G�T09�ce��##Y���w�0�����(UU JJ)WX��M�,!+`%���tpp_-�WVV�PET�Qۅ�m��ǃT���$6c3����������p;�Dqu��d�6����7�t��e�!�)�yR
�� ���w�	4*�Z�Hj��c��L���:��,O5`��k���&��%������?�F%+��A2v�H��@������ X9�!���|���B���W�,F ��n��l�<����{���\�fA�`����H������� �%%!��/$�Ӯ���Q`�L8�������� ���:Qn(C�Ƭ��!���S-;���:8�Y|迒�R�r������$ѩ�^�%%H�--�@���<�� ��:AM�ZE�B��/-��ak��@!W#�s�! g����,��t� ��"<|�W��X�ٵ9�\�1���z�g����w�P�XuO��^p��!RW�577�L�����% d�LJ��8T�s<`���N�~~B��{n���N��*T��ݡr��\������-��_�
�׫��f&{C>ϴ?m���T6Ҍ���V�O�D�u4�W��k����ߡ�b����
�l��2�(}�
Ppǚ�MML2�ʖ ����4|"#Q�s��[�<�vF)�&�u�ǜx�G�����J�4^	�bv�	�ObP ���ۋt�74,TA��s���.�l�����8
�eO�����ܪNbXKmmm'6OdB��O�M��~�)��f��-�k �W���4��� F�sbC�������������Y��������7���5=	Z���͕�u� Vƣ+7��rPm�)xo���޽�)N�<CF^�d������HE��0��f�'Ibœ�V�e��o&B�=�����N"�74�� �̈��u�S}C�Ls�<S������ ��t_���g�^���J���	'_&UHH����/���Y�� 3�:w�Āù�;���\�	^^&�����	M�Bӫ�����,-\������@O��i�pv;�I���=�p`lL�r��V]����1�J����\��lFH��3&Y+�o�;�dbfֽxz���_2� ����927 ���/_PQQ?������#��L_����K �y�'��'=��,,,���
�8b_7�T�^�O��E��@f����S-)_�Y=&�� m���:�a�Y�\̕��ˤ-����?H{��'ږ��AAMo�l�hE�<�W����1ߕ6� ^Ik7��i�T��.rZZ� nh���_S�����G�0Qb#/+0�&Bp�I�(q�;-�h!We�O�'5��s��o�)�:�Xu5; ^m�mx{�ef��!i�I���s�v5T�4�`���V��O�}i�_œl@����F�Do��=��;C�ͺA���Ê:W��1���,�M���j5�Vr��gJ�u}%�� b�Zm�fz>�5פ5�J�>`H���q�����;:D�5�s����>\#�.�->��C��!2t�5pp�Y��H�~H��k�|O]uU��[��/���k6�M[��a��gȽ�{I�4?�E�����ƀ@]s�����[�1C\�G����ԃ�oj��d\bdL�[�+�O
����BҺ7��cD�d�Cױ�PPU1�SKL46��.zA�$��Eဗ0qs+��q�X�,et]r,ʁJ`2_@j��p��J5�G@��;�/�� �"x:C���Yk���~������C�w{�����z���B��8��@�E�K�d���.�c%WE;o��~{��qjl���ؿ���9aJ��pӦ&�o'���
%_�s��=�?r�~S�TAQQr�ٿ���i�d��@�=V�����}|����JJD��E�i|���-�=\j��)x�ŭx��	����~CV6���(Ԝ��d.�Јc%���5Ĳ�����ד� ���	� ��5V��[��n��3�����*���w�UV?�8�3� �*@���p Ȝ���Wn�������$2�@�ǟ�mܑ�SQ����M�C�l�Z�v5�_�C�*�~qj�zK�phL �Q������6Km����;��Ƨ�$?�l�����cۗ�
�F��4w�����{��!�M�<rAAJ:�ܘ� �~�H��q�EdT��;J��iw�z�@�$&"�!�[y��r��l-F�5��+��Z��\pU����5>c��'Ԛw-��3�B�����|pɃ�yKI	"��z����6���|����P}�q	��%�n��+��C|~�Ʀĵ�37��.���k0	X�W�IRon�o���#N�rdO�h;�OM�b���-Hf0 ��%&�t�w-6��v��"�z�L]��������T.<��
�r�n���h\RTR�	�.��a	�ζ����^��A����%����Z/$wfY,�U��P$%UI&&oh�%��Dgwv�F?�[�vD֍�УD<��[�_==	J�,��_N~�hV�g�v�ᗟ&�S᷿��!W�Q�2ȐX3~�ծ��ж�p��*�p\��3�� �*#��=t��@��Ì	]�xkI��ys�
��ܼ���<0��R{[�A >��)+G ���E�7�?&�[C>�S�m�֏����]%���Z�[L8����S��{����������Yk���^IqJM�&%�Jn��/��.uZ6�p]���p���])Ho�5p@��<��J*@����:7?�ݜ�]NUQ�Z������Xn��_"����㛄$��U�|���Z���p��`�����#�G߹����'�e)~�f������4�qg�bhƷ|8 q�����a��sp����QY�q*�/R.6EVUn�?lܡ-�۞$x���˛��r8 ���Y���!C�m�ë#gP�|ה�!���l��׵�~��c.�º@���0� �D�bO@1��D����+6���4��ݮlS�QWT6��W`��Kj	��o�<��9RO���5�Ҍ��=j_����fM���+�+�����9�btm��付;$�`ܰ���$��Sܥ���%dI�+��� 4�U�Kl7�V�.P)�)�����? �����W���T�4JL�tޟa"�'�@�l�-]Bf��at�[�y�WL.���^���tl@�Ο����:$��XTʹ�E���j���ܷ(j���da��#��\����'b{笑��B�2�h��P�T��9h)T��]�;0R����4"N�n�eA�]˂&���Iv���V��E�;���4��s;=4]l�/�Z�:�6EOȵj�~���[^��JS]��b V�9Ml�S�[t	�.@���y�����tt���u�z"$�~p���?/�����z���v]v`O����Ŷ-)2��R��@ǭ펉Vرa�z�n$�����n;�wE�P�p�bf�2ف�G�?��~:��5)���[S]��Q1)��_^&�X�&����U���m�466��2��m?��2����#�w�2a~p���7ɽ����Ῑ��<�.�66�Z�^�5�Bχ�&$1XAJJJ�@Wa���c�Sx]F6�]�p��������Ɨ�q��#�űGL�k)��D�W�;�=�����4"�Z$����*$��o�z�GD�R+��\�(a�^�4R,�.S�S�~%�|�o.Z���j���r(F�����>F$�Y�죄?~��nJ�V:�R�u����9E�	q^��x�%���[Y�I���!�ם���J�1~{�s��b�����Y��_7x��8��M��\	,�b}����U7�Q2(�S���/��w'�&+��7Aa䛂^`&�K:�O��F�5`��%Y�<��l�c�z�e����(3�c�+���֨,�NY��.��c
?g�ܽχ�oꄆa����=\ 2A���{j��E�"�A �)�YZ��E�X gP�} �]|Y��Q�,�M�5T�Us:(��a����?������Y�pE;�A�E�˟��N��o�'G�j��RMy�]/����ٱ���ԥ����
(i@/��8K��v\ͼ�B�YѺX8π-��f�O!�A��y��y��������m��ǧo_EXL��6u�(���z�������]�Уc��W���ʯ�S�{[��v�ـ�<�g�ui)���������:�|DSw�i���aL,n_j݁�I���N�b�e��Sb�c����v�OӺ�O��G����~��;<|���'<�d��ҷ�[���CanŮ��3O˃E�����vB� �
�QH^10��F~%s�i�>n�Z�=p��k%Z�C{�z���
& ��jA10�p�f�� ��W��]��o� g��J�dh�.t�=vh��`KM^����ɭd>�a����:,� ���M�x	A�4-+wI���W�j���[Xu��|S�쬔�`3��8���	���%�de���5^�J�?d���:"7g9���bM��ͷf�M�ĺ�*D�[q C9r��X��b���s��a��1��PU)���^Tll�eIT�_�o{���?|#$}�R%mo��3m��QK �Ű�i��IR�>���V/�"�@�g��|�5.�w�>�\]eV6�*�u��!,\�k\�!��7��*u�{���4� NZ&c�^`=릻q��~��y�<��v�*Ev'J���wu����� Ẑ6`5����=�������qv
خv!�ħqآ��M�s��LG3#q���7	���7�;yzܔ腪�7�ւ�ɘ�oܴ��������xۮ��¥n2H�x�D���Jpp��2/�)D)�4Xf�:���orM�=3^���I�56��ğ��ZV=��l��矗*"�]M_Y��x�Ԭ���H�}��F�u6����
NNN�Mbdh����MM�Х��W�����}�ݡrE�}菗��s�A�X�E��P��o�]+�(���]RUiŜD8w��Ŭ�R�p� 
�%W�ZZc�]]]�e�ȄWH"��t�#|Y�W�ٹ:FggC6��s`�&�-|��O]`����g<��`���7�[t#��p�v���-���O�h[{�3��(�\��Cm��!�T� Xԕd�i_Pu�.��Y����n:l�k�|��I m3iQ➏�,����@����� Q�J��Ѩ	��)~��))2^.V��-;���a��曦�:y��xkn�&�Ԁ���� w:�mR�a�|z��t,쨁����ɀ����{G��f(5�^��N��~�ӱ\v���%sXd����b������-���Vz,�{R���~s�UF����4�pv�bpK�/X�y���WD���( ^'6��oJH���BU��\�KYDY3m�� ��T�b��sm�[mP�<`N�'��K��ոs�!5�@���9�@��k�<j���;Y����2ܗ/_��jF5�뜎Ib:�C�xп΅���Kߜm]~:�l�������Hv�QTYfA����4��|���t�o;�����y{���;".'���}/����߈�oY��n���U�A��
e5s���٬ac�I�������������Y�Y!���J�\�·� �U��C�J�����JD��-u3�(d6�ΆOH˜�뇯�G5]���0ķ7��e7���a�! #g�8-�)ض�v�C`�i@�#^��C~.�	��Q�����_������C7<����W�o�y������(d4�M!C�N���7�)L5�g�NLT���gz�Yŕ��\=K�M�9M��S�`vv>HQ(�o{w7d/�f����B�Ҭ����\�Z��E5i���^7`L[yzd"���`![ݸ��^�O�>|�����9�{T��9X6�۠FMR>��
g
���_g��s�iݞ�g�T�庐�zz�o]�H����ʔ(��̴ܺ��w�777�eE���*�{FGџ*��Xk�%j>hA�W�UM��.�p�s3tÁ������f|<<��>5�_}Tp���gG����-� ��=��w~c$�����o###�*�S����F�ۃX[!Y5WŎ�ED�S��w���|o�_�s�m�,�Z��E��h�La���5xy7_���8������M�G9^�vʿ\۩9��#�w��X6*�Y#(��������ȅ�?W������T~^��&��X�3��ړ�w�Ϗ���5�����Չ�GP����{�{��e~��=�vV�%%'�i��h�q�L�XPXU��=��Brr�$$$�e�!�0���^\��쌫<j��T�<�~���
e1C�A��X[���0����E�$G�˫��@���628Ԏ8�.k�R%fdD�ï��]���n@}��c?��s&E�>�wt�W�Ku31)��\ᑗ������Ĭ��}Ee��ؘ�\���V�y�)Nvtv&������	%%f,�Ħ+.�;?( �#-L󷽱���B�/���"����7`ͪ��G�R*��$�Z�P�͛7C�aFf.��i�U���̭�<�` ������q���J�;E"��>��4K�Υ��##f�X��������}0k����Dx����i:�l�Aȓ����H�md������(o��qM:o�ǛW��I�����:����ޖ���Gkȫ��j�tt�ΌP�*�h<�I�.�㭇��(�zP�Nv?v{-\4>�b�X���'����B$����g ���m��m?��($�:�-���ҝ������ry qw\��?��϶G+����VWV�C< �����.w��o ���EEUX��5`�TB{��X�e���̼1[�l��f��iB&�������p�5660+r�no~3��d@�j�^��Jg�[lN�_z��ٙZ���f����IE=�������Y�wQ׆X�gȫ�@Mr���rt7 �P_�{6S�t��w�U�NC�|9����"� @	�J�lğLm� �w{mԢ�Z#+�ub"���[:_�<i�/&Q�>�7�=:�к����Εw� ͓/���AZtTN��Su�>kТ(�E_�|�R�r;m����Y1������''�O��+t�39�oҏ;t�����;^\�gj���P��oh6`��o��ݩ�7��b�������͟K���Ύ!���S�8Á�Y����O�X�*�X����ʥ�<yh���4*&E�zcc�oϬ�pc���3��g��[Q�����\�~
��<�ma!�ǈ���l~g���f$�OY��`�c�@}ϛ�U�1�L��]�����������::.'?����r��Y�y�.;KA�.�H_�ST���[���I'�yD������]8�N��Z�k^�z�p�C�D��a�)d*�z2��]��[3!1�u�;|��OG��Oٚ��G���Ց���ӝ��p���J�8zRi��:/ �R��ZjKK'�,�pSu��R�U8��=�7,�A!�n�h��NЄ���aC֕_��bx��=DI���9���I�i3�C�,�����{�ʷ[�N�(Y[�:qRӰ�7��l������X:���Ǎ	�f���(��;*�� �s��;����nX�qv��mii)�_e�8'Ȩ Ȥr�ut@Ъ��=��ʹ�O�s���&��'��a�Jc��<��Br?�GF�}��Q�������OA�_k�{>q_�~���E���k��:������~L����h]z�|���S4a�vLd6��������O���Фn�cm�#��(��ɞ�g��I/�u�Ј�A��/�o���-J�ż��b�8T�����f6��i̚�X��o�`^1S�<y���",hSEL2kj8:t��헗�Ar2E7i��kP�[� ;��R�~eո'1��"^OA���@lr_��t,晳��ҍ+���^@̾�  b�3<_��]LW�>m�6-Y�M�[[Ce#++F�Ƕ���b��Syp�ug�
�%�=�x�ֽ�*�R��i"3�c�fryu��$�i&�{��U*��Ll��+���	�����t�:��x9̳� o���oW�g�6�SՄ�����.Y��Uק�������O:`E�Ĉ��I�A��Lx;�-�(��k���Q��s�	��Ɋ¬D�0t��
-(2����{x�e��|��wQ���rq�.P���۠��(��C��999rI��tBc'뜮�����`�yo=������dtuIbLv�*��L�`�h-(�N����p�QN�j�ݱI��4��T�x�hվ��_�����}�ɍ�$������3�e��i�M}��̗�A�Wܣ0�Г��<�KeSP+��|`�Jـ�ݧ���_1�j1!x�����a��Y ��À[�X��F]ഉ9��J}�Pt��ixr�_P�~��+�� u_�
i#s��w��%����s�`�[?�������\,��>�2��1*�Fmb���]�#�8�l��k3��|��I�ҹP�qt��ΫSjAߢ��L��MQ?�n��9X;���8v���N4�hW���w�"i�M0Wqƌ���)�qq��@@A�H�i�c2U �͆Y)�?::�y�]�9�R헞��2����H��(dY���7Ϥ�/xsI���?��ɡ�.0�N,��?Wp�d�:��42.vܛ&p.�[<��@��})j�[!P��~Ɩ��Q�q�@�P�y�a."�3�c�K�����-b��b��'s�ltK�C��s���l��͒��7pA��M� ���~��d����^%f��w5��t�1W�'G�4dR�0ͯ���e�lZqJ
�H�o߾��ȵ���O�?9�֤�^ߝ�{~��DI��#�:��cf�4\?�*���ɞr��b��r�c�-;h���g ���@E*�T��cS���� _��U���&��7���,�2�S��ZXh��x�?|?QzCNHb���G۾h0����H������1��?d5g.�7���F�?���Q��w*�or�|���{�/��z���\(֧�NӇ�O����o;�f�I�c�ݶ�rЫ_$>�:��B��Ю���R�0�>������|�R~1i�v��������tH]�S���t7"\J�����A���C�I�������{����眽�^{�3w���e����-8��8��_�C�F�X��m��˰W�w3w��Jڪ��z`8��͵��G�šV.���Jc��xm"ȿ'�~B��!E-�"jk����W��+�5�D������*��y�P
���1����H@+�H�m[����!uS?B��?_�tp0��Pڅ ��d�Y����{H����,1;�oµ
h�A���-���t���1YR��,��g�e}"=��<����>=����^@���d��DW�2J��-�}�����\�o���e�`�����N[ƽ�\N�R�_D2&���3͹Έ�Ӳ�|�������MRi���\�z2�e��(�F�B�?���FTyT�n�삤��0�����2�JB#_ ���v��nߟ�{���ÝA�Ÿg����;:�����/�`R�����W��U ��[.���I��`�tŰ'�s3��[����n!��}~�V%����O3ޖ>)�����C}?��B��q8߻�C�{�%��Dq$֍��Zy�b�w��A���arO�Ӫ���eM����76�����h�vv�\�)��ȼN��%X���2�*Ex�c{�@���
ew�Aw�UdG�"�Q^I�2��b�e=3#CFAa��l��]�g�Y���[��{&��s��:�h��:J2	=�xU���vS"��껟j�6���N~�?�Sr��k�e-ә.e�s��&h6��i��%�k8���8��E�Q\R|X�[�˴z���;�*�������A��;���S�j��F��&z�,)a��j1	� 1�\ZZ�	4�#� �`�xP�}|s�&q?9�uP%����ۙ#�����=�i��"k�j�DG;)S�F��ӽF�������)N�������'!l��nBOu��3Js�?$����%��i%���X(E���ZVK�x�t�r�752;�0�ۤG���|t͞/�zs���kx�M��ƖB���+m�8�>V�;�%!1��~vc��U�U��ێ�[n���I����T�t���?�M�*)\G�	�o
3c�h���84aR��ʌ�wR�dw����>	{�%��X��������e��z���[u���.J��W2�s!6R��@�1i�	��)��*i�q������j��d:�.�$�1Յ�5�x�"Ump,�w��y������`ҌA��բ��6z����� �H�Y��[�s�F'���B����T@� ��~�l��oV�C�u��Q7k��q�vtd�G@�ՙ�ݲH��/acS��Ч>�]_b�N-���0�e�$���*�>\�gʻ�i�Wv�HJ4��3��WGHuc��u`N��w��}BҼ���c|-�ૅKG�U�+�D�A�I,�����)8�hl)e?g�E�zη`���	�3NU'gfz��2��O�3k��b�5Wk�w�J������L�t���D�S���%R���0p�TU�~f���&����@��%)kF���/m�xoŏv�g����}E�׊�A}R)���W�9���:˃Gw����9X˚i�Z�ݐ=?xِ=�K���Ԯ9.��E̹��jg���.<��������r*�럟[?����&&T��fԙ5h���qxa��ז�^�V=I
Rƴ-�g�0�����E������.�{q�5@�5�fw�m��0��Y؋ &���X��bI��6^����n���ꭒ����j+2&Y�Y� ���4�������m��`b�{�=��_H��fz]^��ݴ>��K��`�[���0c��Y���mo��E���u�{qZ��*���O8�:����?ma��B;�1�^�!�T�pE��c�G��t�k7�F��Z����`�+-��~%����Y|���^Q���O:VVŽs��C�fwLr!�۔�����o3�(��rZ��p��ۺՌAfuֺA��z���i
7 +a Z4+�H`���^��c-=�7Wa9mw�B����U�=�e�+ã��W�u�#�O��W�n~�������"GIgZ_�D�t�<F�9��}'ݤz2�۲��a�Κ?yT�A�M��jdD���RN�fl�%!R���<�P���
�]�!i�c�l�	����U��T��5�v>�V�R�)�5#F�}���N������@m9������r��^�`�[�9"W����c�lq%y,ںɭ]�ޟ6��s��e�2-�'7̍��#�Y�ZB��;Ы�6��M7׾ �|�b�W������j]�ܘ�H>t��
9��E*c����f�r��2^�N�t����g�O�D��yK�V�����t�`����ի���'�4iiy�K�Zs���;
Y��N�������j�IK�����N�^�{� &Z�BSSSe�{�W��?U:G�s�U
��/]Yt���l��ܯhӳuԋgÖ��:9q���+��l��\1�:W���z�x�}��* �?�}Ê��6��#�����4�{�Ib�1f���2���X!�X���Ցdg҄ԩںS*�MǟD��4�w	�xQQQ,,]ק�
��#l>tCy��L�-�$�upbۣ���F���wĪ}��}n��tEs�ŭ���0i���?�vSW�t�D�<{#l�W�c!��{�_p���<��M�5A|ʷ�����(R�7��bBX#�+p�M���y�lu_���±*�V�aҧƾ#}�I�-+GnȼY�L��zWU�g����?.���Q>Xh���pZ����}��uܥc`f��{#���4t|:t�k�ɟ�=�����^�C��4a��K7��bݖ�A�v��t�U{��r�wqz �X�$�A�<�F����ܖ��sunl#����\Q�� ��;��a���|���H���پ�$q2���6��X�����
*��\Kk	qq�%v,g���0��>�CO��4�lg��7�~��ѩ3�>��pd��i�xT4���k()��p��Qځ���Ԙ������h�i��cH�&L4���h�R�H�Ѵе�����L����s?^�[����xt
���O��4b0n`[�ޔ��B������B�U���/5�Yn!�'d�=���7L�ӆ�����v�Nb�J"ߛ����}���e8�{<��Z; �0�8 �{��j�� 6�����[éa�<�i7ϐ��M�`i�:ðև�� ːL�S�����<���e��R/447i�
�E菕�u}��|��h���Q��H��`b?�*��
G;aO<R^뮡��l�pl��G�Q~�%2 d��&�AU��e:�?���/�º�́6�MM���坓�C	�	�]����j�]���M,r��z5��.
��Fv�i<�mЫ�joP�#�ON��'��:]wpxD�^�}N�z��)yT�jE_��j��G�(�4BÑ���>��x�T�3Ģ��T0v#�;]=Q���_�x&����4&������%�D8:�.2y��Q<����_���Q�����}���a�#+�/�?�+Gl���u6<������jƸ[�ylf���8�+�w��jj�&z�Jz�Ovx����bE��t��Nt�cw�$�������9~��E��b��F{����;� �\.��3�+�% d��ȍ��]|�h��w�&K�7|��H2�����"���*}�)���t��;�֫%��:6ߩ���j��{D��E7N��.Ӧz=(�H�UUq9l�<{�Z?"=!�[|y��
 Lnv�[/6r��../����6��B�!��.[�bOa(�Q��fR���t�[���ᮙ�&��_��g�?���3Y�J��v����c�<��\��}6��P�V����Q{W��^A�X�����pg�kH���P��(KZ+̡�!1����b�C�F� r�sǫ��]J�������Յ~o$\Gv��8J�����=LJ�����}�{-��Aȕ�K�\��؜����@����GbN�\�}k6������a&��C���,J�`��%)IIɁ������cIU3$�0]����(�w/D
�U��l>�Xݦ{�h;;���e�k}$5=alP�?2ש�lܷ?�������J�����Pq�F|����-����6<l�N�jAF���	��6@)�9�ܶ���߃��{�7Ʈ�1�~��?7?-;o2E�C��_?5P�%�%v�_^;m+^\8��|$~��Ș�N��_��=@0�K��J�V��<�����4�:
ማ�-���d��4�.�H+�%�:_�*����(a�  f�+C0T��侊Q�]��gw�n��;y�W�<��@)�MԴ�ɼYN�Q������;N>��t��f+ō�7ɱ�ha��vS?j��`_gD�����l��f6�����}��"@�6�f�7x�n���.H���kZ\�w>ę������$���h*���o.V�i��GL9nU�@���O��P[�cn��e=)@j�[ւ��Uf�r�"W3��P3��9��hf}��5����A0_HH9|���������+�%|��УG���K�C&�Mb� �#��#c>=�3��{�NԨ�j��<���púh�:j�O[N揩K���.6a����*c~�3w^^^����o�^����|��O*�� �_6�vm�x�3/�I�����s��mQN���/���㼼�y���T4���>6%��&͔��C(�Մ+�5X�^!UVS?]�uC#D��2�)������ē�^#�1����t7�՚�x�7��ps"�ɋ��p'�����1d��g�N��������9���R.T��,�0e�t8��7r��藟N���:K،��y>G29E��Vk7�N�sv]�L�8�L����b��TGh�:�I%��
��q���Nh��_`��"DY�(++G��j϶��Ul�u�]�ox�N�������������AUm����B�P�XN��2{��K�n�dx?���eK+�N@#�O��/֮��r�X��	��9����ڼ� O6i���`c����2@�^�8���H����y O*�g0w�@�m�v�Q�a�%�D{hF�^c����;H	V�A�*�Y"n&���tA׹��]���Z��W�����6�ׇyݲE>� T�FQ�{��4펊f�(����M�Я_��%��^��e�RR��������R�-��������2v+׵rOޒe!%�n��ނW#YZ���'^H�(�I���}%_�=�]��%��㝝���5|�C��**�'�l��/)��k���X���`6���2o�ɷ�[�6�,$�2�������}W0*.DK�����$O�֣c��ٖR���&ڢy6�\L��~�m�م[~�������%%�����6s��pW[[f�L,������Н
f�4���\��?4��6/���_t+��3��W����B3ݜ=�ʞ��l�L',0�:�h���'K�B�fA�ϊE=/j�EhU���O�l��[�@����ܿ�~Z�<E �U툦��q���͍w�L/�sD��k��YH�^F��h�7m�Ƙ~�?�F�P��z��q>�k��t��Q�c
�P��*Q��5��~���W	vx��O��Y�67GކzN��!c?���-,X���oښ�ZT��O8w���3��Yc��qxxx�ƉЬ�H{X�֨������䒿�=�Y�_n�<��:<=�K�.���T\�۾ɌM���'�HG��f!��lH,��T�������é`���`�/0S�C��$ ��6�:mPH�1��x8+w3[���@	�8� �Zկo���4}N���;���k�ԍ��ֆ��	�,V!S�3������7h�@��&��/���t4̵��@�@�|�w�I	��l�[a`����ˍ�dk�#
���(��;f�� �����y�xˢ_�r|�ջ6� ��W�#�i����ۡ��tv����X� /�(R�e�jA��~�Ύ�=��E�W�qPӯF2�L���ʜ:.�k,�|������=�.wLjɫ�zՒ4�/��a�Y`�RQW���/8�}��3�T�W6^]\[Y��潖,& ��B�bt
o�*���xxys[��t")�8�7��b��c�닏�5�j� �s�*��lSe>C�'����iűi�@�Z����-l�M;����)� Û��f+|(���4��u!5��γ\�<��yW��ϻ�/��: �2��z��Yt��?,WS�%^�fy������@%?ر�J	Zw�2���G�#"�u��b�p�5�T 1U��/�����jlߞ�,��~,����x~���qJ��n�p���7�o{>�^��
,ыX�ӆTV���s'�$4@�b�u̪��XFOo1�+==]��۵�4l�<Dh�|Ȫ�iõ9�.�n�3�t�\�Ю��zW9����؈C��ȓ�<β�<�R���5EXYm)��OO��^���4�?6���>��o�rp�3"�U��c��\C��`(5*���JA��+��M�N[#�k����䘞u�N��`�u��.븰}[����e��Nm�;��_�������m�����z�I:_�� 2������Đ�b�#?7�=R�{>��j�ב��I�����e;@�3���%G�&a6��.��&�8��r����{$������י~���]�W���ɺ�Z���t�
%�%������a��8��ä�����3��}H�i)���i��� �4��D �n7___��Tb�*��~�.����=%Q����ϔ��?���%�4[�ٱ%��" �0����t�,�ֳ�C\ݪ�,������U�l����O�NJ�2k�����p���.ߩ��{�RBK��'] ���[�ڏEՐ6h�~'���֖�p4��4볩�w�*�|h�՜݊P꫿���r�p���~ш�rx{󍅈�l����%[����KKK�Q��ƀZS�Դ��ef��X1O��HJÜ�l(Vo||):�Ѻ�����}�\e���D�����ѳ�[���%��#ݣ|����q��6��
$�	����Z��Be"^۴]�4�@=����x�	��߱j������	 �����l�#�m�C�q����xc����H}����j��U_��v�+-�Sa����H��q��&�����;��g��a�k�WO<�Xm݇2@p��*��O �?�t�
�
�����`Ij�څ�?��8P�/&��V�Z���}w��w�j��� ��S�
�S����Pf[D�'͢�
ˋ�#�<���q����^�䉫�>�����l��/�;o��x϶�fx���0;��Cѝ4Sgh��	�߻T[�:E��b��z���WA��J����Gxi�K0�}Ǣ_��e�f���RG|����n�jOTgn�����*��L��W3���,���ƦW��M��j6Hm�������v���k?�{\}�S��^�����1-��1���srhX��Q��5�"H��1X =YpE�(X�;��뷨��/s0U�F�7����S��l0��F�������h� /]�לoQ
��|w��pL窽��̲�p��#��;ѻ]��*�w�k�]�c'	�hP�K�n(3�_����#F�e�q�%9����'uzUsY���Vi�Q�ّϳ��k8\����Ϻ�/KW����G��9�[u��jC�����7��*s�G`�S_/�1��p���qD߫ۘ����|�ǋgW�G�|#)�V��"��ټ=9qR�	)�s*j(�(v��$���.�|���C&��U���<����S:�J��b� b����5�;DV����e5;x�]�}~r�Yk�-�2���g'p�a�GF"n6h�u��q<��\f3����.d�� �(�����!�V�{�k�P�h� �7���'�g�����U��-^[++��'�y7���0��3�N1��TAt�Ej؄���"(eR(���8���dB_�0�#3'.���T�s�a�ߴ��X�x�:92u�:\��[��yT� y`P0��D�#W ��ۡ��2YV��^�𲖪c�a���C�
�}��XÕ���#��U��������(�i
R���?���6����6W�.'��ȁY�~��*�_��$������o�m��M+0QH.�9�${�p�� �,kw�D:8�"�
ׂg��Қ8��t��#��nu�K�	_1R	��`���!�&��4��������z�u��r��%
�%F�V��&�	����[����\zA������g�F����:s��=$��*�-q#/�S�)���m�mR8x�ܗ��a1=�+�^�!�6-�p
Z8ȝ����Ht��˧�N���2�l������q2u	8���e���{��R4�	0��B�EA ���'i`q4����Ӧ��Wi������7�2�t��zڠK� u�3�2�0g�FtP:H�2����ߣ����w�IiD�	h5�d�E�Y#��FQ�O� 3�ƿI�<3��i�pl͉rO,���l(©�F֝�z����u���������g(}��H�	�B1|T.GC�ޘV�s$��e�a�+���w�4��ظ�v��/��ϭ^1�9eD�Mx��7ެ��G,�EjB��|r��H� \�Ϻ�����j:��܍M����>��7���(n��/�l�a��s��1u�Y��\��`~��뷃�O��#A��Β�%����5^qi�ɺZ(ziۄ�~��C�SR�^����U�\��I��<pK)��A������O�
J�[�j_����o�O���?��8,�5@��b�������0�7���0���>MT׼��hg�m��rB�Ѫ�4���|E]�8�0�y���	�d���A��(<]m(>^�3F?$	*N^<���NVE������bJ�:��B[$��ğ�G�K� I�Q]�@lo���~QL�p��K��=M�&$l�Y�z]0���k�RJ���� |k~B�x�� �y��C�Ba�Op���h$�_Lt�t������(]>mdb�	�w	c��DȂ@����]K �WP},U���������t��l��P� ����%�6	�X��i]�>�e$H�T�CQ�h_�ˡ�����[+ex:��,��kq��#�tE+v���z~le��'>�A�-{���C��n�I�D�<�`K(v��k��͸��隓%VW�0(��
���'�-�ɴ��oّY���*��9ZA�z#`O�VG(��}$5��!5�~�'�+j@�-,����v���Q׶�:J�>�Bm�#�^1���Ԛӑ*n��-U�emw+*ċ�l��L)�bE�>�.^P۶y2@��;8�֏'���&��sד�Eߩ�O���d�5�t@��~�B%XZ�pӆ��?��vRQ�5��(��:���U�8J�x+v�O[h����V�:�"��[�ˣ�3#b�P�+.4!~n��xt���CP��,A&.�ʥUZ8c�|j�h�~l@>o���W�"�a�
|�&@��0RG�Li�l;\+��;�[���z��Ci��e��5�Ƹ�N�/WdX(�L�l�Bw��f���=�m���Q'�h��Lp>���;����z���4��զ)�SG�êv�x2CY�*��w�P���QG���\��ty��u*�7�s�;�O����U�/J�0(���������G��9�WO�D��.�H2����u�v��0�r�@,�u�{f�4�O�w-U���y ��zy�{&h�n���j���k�{$�5NT7Nkh��4��5�WETt����P��yr�7�
����3]M��%���󮫴7�L�ғ������H���ۻ���"�V�l���J3�v(��&���"��q
����n��7"��-����l��O���V�����GrhBYKŨ٩�����4TF��^ �iB���+ili�`��ͮ���H~�Z�VBqpY�I�u� nV4�XSlG$L��3���;ݮ���H��܊H�J5P3��?�"���Kt�`BF�
3!�߂�搋�3Apvm��L����)l��J	��)
C2a[�J�h�Xa�|J�Ǳ"�?@��YΦ�[�|��M�̳4�G\�s�����@���zz1p��U���Ԧ(V�-��;*��F�*�y���z=�@<}�����ƙ�!T-�v�j�� A�i�&�w�8��.�ʦ�@���N}hZ���`�`2��I0��5�Q��#�`�X�p4�� ѷ2>G�	?ƅD���T��0y����=~S��+�n;�m����j��^ )r��r'[�'W�Z�%����4��m�"n��%$
X�� Hgd��x�\�Ƹ5'CO�U�n�"����.���)�YKGUq�!�@0����8��YWK��#���4�	=�����NK��s�:����� �"e.g
���LYL��JT���O@���vGV,���{��W�w���TGM�5��o��п�Z.���2cYV�!g9(���G1���Lԣ�T]�q`��L@"Y���P#�}��G��=�]>彣���l5"�I't�PZ�ٯ���ƽ�$o�I�o.�JH�?�<�&���yqw-����ÿ�'�}�E9��~�5�g�U����_�smv<W+,m+l�5RW����`Z{��qkT ӓ4�es��#�y�VF�do��b/���ۋ£��\][��=lW�U�b F��"R\d�'�5A���	V�j���ܱs��+��]����3�o�BJ�)�mI\�:\�&˹��;�-w] Ê�'&p��ـ1 U������	�T"���Ԭ�2��>t�;�@��#̛^���{��LD�2P��_���P�����Wv��J��A�,���d�4��u`��a ��Y;벽�~�@�����l_��9�.���x@t@M���f��X.�$����~�'���A*z(㣒��e/��K�Z������%�eW�B�����>��4� ���6���E�	����P�4$�.Y��z.��;ѻ1,���膉�e��~�#���\�E��'s�d���=}�OX� �lAWq�˻l�a�.��G��!�a�؋q��W��c��6jq���b���#��b���_� 1�l?DJ3��xR�f�4J���v	��Ct:�['3���[=n8UHf��e�5�V��'Ҽ��4j�'R�^�Z���ȉ�YI�Y�HD�=��$r��b���բN�}��T7f[9��= q��t@�!k��}�U���^�����S�5�Ǯ�0h�������k�k�`�@<=�xQ��0��ƶ�l]�Ȗ�e��i0@d�n����z3*j�x��= Lv�L�����D����}}w�` �ˠ��0���.�P�./�a�(/��(Dۛ8��_ ��+4Y���w���0�^����*�X���VׅZ!�[e���JXe�`���
i2z��j3ļ?��k;&V��h�	��Z.J�{�����z��#a��E�YI�0�pXc�~��c|RF��݂T��f�5�sr��,�GB�Ǐ\�Z���Բ��}e1g�3,[��*w'�EE4X����Vb�Ezh�Î#�ߛ��h�����p��"�x���B(�ZV*k�Á��HGܖ���,�HC
�-|g�}���ۿ'Uh���䭸�3@�m�N�)�JC��%A��"�����]n��UELL��(�H6x�'�3�Ą`��>j��<��%����wC� ŭ�ItA �2�R;֍�0���A �n���N�00���Oݓ���oL�����'IJcM�W��f �D��Y�����v}�Zw��4ZS��(��F%i���uXR��/-a'ט9�0�Q -H����G����<�
sL�W4���UV2sR�R���<���j�!�R�d{U�jt�}���>���JM�k�ǐ�Y���uW�� L���M����!磡//�."瑁���
�K���Uv$J�0�*6���y��y��(�?%��q�/aD�O�y,eW����{�P-�� %��� *����(-�{K	2��/6���L
7$K�̵_�#<� ��"��Ֆ�t$��+~!�Wt>��r��\ja)f'P�C�ӀN�bT�	[��D�0�3&���5�����V�f��Gx�6B�5�)+[��g����?���c�£��.a!�`c�#��Ϝ��d�b?����j`������^���/	�^p�&�
��>0j���M9򜗘��� �a�o��������}	�ʔ����%�p���D����7�ŏq[��-�()�Y�|@��Xh�d�-��u=,�'-N�#�B��@%eE͈G�:�s�p3pb��9���L��|��{2y�Cb]^��'����	�|me<���i�������#a :8W�����w�_��u$|�f#�>�y0�s�(�9��;�H�d���y�����f�=)�����\_�,e���Z�@��NX�_�<�r�l`)x�Q�k���1ZҀ7�#����B.Ed)bp��B�]��%�(���yK�6}��/�o��m`д&O_maqm�l�����-�)�⵴3�����T�<��:���5�8���V�b�4(O��8s{)p�.^�E/$:�0T�Ƌ�����}!�#��ER\�p���vऀmʐ�J�ԋW�H����c��Ivpz�7.j�)�4��;nl����<#ۧ:B���O��/�|�&��A��NS4����׾����*��5��ߣ@�ZU���3�;�[8�c�}�V,���R�|	M����U��[��0@h|��}#�>E-���'R0��=�CI<.����[� ��|y��e~p&�nz=�Ǉ�����C�>0�����ۊf�.B��x��n�l�侹t���q���,7=F���ק��� ̰��m  d�|ݲ����%����z{fE3 9Lsx煘��������v�*��˨ ��<�7�>�C&nՁ5� ar�@(��a�Q�K��G�k��<����#�%P�Q���}i���#����ca���������%\���r����\O�b�6�󻷵3a^��EV?[@���J �#ܞ�0�B��a�(�(Q��n`m�Wwԯq��ل(b�&
	`c��(._����8t��`/~��m��1\&wg"0��3��͍}Û4�"�J��U��Xʱ�4u���8Y�vCP�l�2�P�&
H�"Y����{��Q��p	[�{��q5Q�(���~���\\\��:w���a���w~/1��	�� NG	�̵�y�J"� 	��K���@v'�?�"��D�J�SL�J���L� 20�vC��X{��a�	�!XOn��{`���8�D���A&���������һu`�;��m� q �����'�4���d�����Q�������#�<�x-t�+j�ut�=�h��37e�]�QT�	u J�������o�f������T(�X6�'r�*�b��}X;�@]�r����]����P�L�j�����}�Ѹ���1��ZQ�c4{ip+uy}:(А=����^�+�����sűa巧B��څ�}�V7ԅ��PO��-�|[)�-���1���YEE�j7F!�䲔��TMX;U�5�g�k�r�[m8γamZv8��Ȅ$��=�_���y�.�`�]����p)��J+�\�a)s;vK@��784����{��e����U���~-5�P��8�p�� R,�#�'}�(9~�=�� �P��`
@�#a?YːܯE�x�[$��{D�i!L]�7ֱ�=KЖB��9�;a~�5BP{=	!L�{]���5��'��S�R)+]�&�L���9�����z�YeJ]EȆѨ��1���Y�p#�ǡ��u\�e�ץ}�7S�|;�H(F�O�%Bô�Ko�Ŵ�mh�R�X�_��d	��tuvu}�p�%��~qy�6[i�@c�9����f;й5���wB3q��7�\�
�t*'K�	�B��"��2�Eӈ]r�RT������}n��E�	�\����36��^�p;ۅ�*Cpm-p�Bɔ�\$��s���X���s��E��&ȁy���5�u��;GG2:::�g�['f*����G=����{������ʍM��O��C322���s�566�MO���H1L-ûL��G���6�m�cT" SЯ�~�ƶ냖_퇱��˱H��An��,Y^�E�y5u: �Y�����:�Ņ��vFQXX���@��}
�e@�Z�1�&X���ż�Џ�� .���Q���#;�47�3�cS�sW�ۉ�;9'�Ϸ�� �@����H�'n϶�9�[��
x�F"@�|������{ֺ��E�A�ք�k�4 G<:�̀v*m����غ���C�RZ8E���MTShэ�$�a�5V�	��i���qX�QummN]/������K_�����|�hp8��Ř�vf�	��|2�H� ��u'���-��Տ�^d@%�1��Z������XYY��e/ܧ�y׽�� �S�}�z��N�f�L�3��COOo���ϝ#�ZX"��~Rm��S.V��u�wH�ߔ<ȼ ��>�9z�j��c��a��9~�f��	�ą������{[M�0ft�_C&  ����W8���=�>�¸�@�oXJu�X1���Kzyyɥ>��k�����daRԛ�ᥐ���[b��/b���U{�� �⬷��?G�5�T��`�q>Т���9;;'S�$�[1�����ȅ�Hihh�*�$��r�ڙx٣�n4�d<�����f���Ǒ����a~����7t�B"����s�&J�@����Z��6땐=?��ԧ�$×(>�z2�U �&:���aU�~%����0l�����M��' 4�����|�?��1��ٗ���~^SP���3/��0���J�@���n;�J�=�+3�:1!��ǫy����|���I
��d��%Y��}�pqq��;�s���}��;�Q�3\��v�{�D_`�ɓ��ܼ��M��rHT'�k�ʍ�\c�������4t`�����6��r��fCt���Ո%�v���2$2I5�8�~%o�����h�f�����vŚSq���~Hq�@�9�i:|͉D�P�[Hʱ|f9ί�̙&�G3/��	�e!%�XL[�KG���i/P/�X��Es�A� ��6Ns�gT��VT�ሜ�l3��BMLg�]z�Ǆq,MWݵ�s�6o�*�HU閼4�-wO <2�bƈ��,�J/.��q��nD�N��,��j��#�Ԓ��EZ�HN4�rĨO�!go�%��y���H%%�6�}˪�"�6�)U�s�k!�@m4��l�A|^ҷ��Aϊ�V����|M|z��K��8�ė�ؓ�j6&�N�mL�LZ�]�h��?<��)~�x���^K�ΐr���`�q�>��+�@m3�|v����\M�̀�b���O�V$B���7���C�kWLQ���$Ԋ`�~j.�!�#֬��Rw��`����衯mVC�G8����oƲ!(@��>w��v�3"<u���0u��F��:?�x��p��R��E q/�3�\�5���˲�~#����P�g�5}����~NL�0I�9Pu�ҫ���e�&$&�����4���LS[@�y�AH�Y�?�p��x�H��ok(Q``�5vs�<�-������ݏ���ٯw��"6�Yg��p� ����aw�\+#�5a��)�6$Fm�g��,m��a5<Q�[@�nC��=l���N$Z����#�
��Խ�{��䵫
��c�����s��H�B|�Z=�bh_�(9�K�3��n0�����im�$�d>s!�IP���9�u+4ǣ�������>c��Y��\	t����[�[���	�c�|p!{,��"|���0���f�@��Ɯ<���\�F�Lf��O�����t蕧�g���2@7�b��z��9>j_�wJ1/"�1;ȼZ%��FSd��1������a��#Ȟ���i37l"jٟ���k�(%*�h�A0ً��`������7�g!�F�s�U�������R/��3
aM����7�p�}���P*�����5����pt o�H]����K�����_cMr�w�{�L,.��v�\?���7��!N�w��)3�rU?D�$6���Ek�q�=��3�V�Lj����tz����B����gl[�D�����-�#�'�3'��F�M7y���] }��w+h��*��Cz�l�ȫ��4��l��V�����`\���-����g���1R4�eB��C����p�N#q�sOpR�� >L-W0ȥ��_:������D����ز_����;���,�
q�t�Gڪ��6�@�g�j�1��|>�A?�.�4#�wk'o
�����=�#؆g�����r#�~�mgƻ�e
C2א�?�$�b�^3����D/�����x��,�{���d�,����L颇��T��p�鏜@"X�fb�U�|�5ݽ6�-��c���BIIik��9�)��W�k�^��W�C	��4v?"��}��7M\��w�Ɨ�2�l��:���+sZq�������ĉ�@���l�Ǹ���ͺ�|.p��w�(�l�Bv�l�!{r�H�Lr8�6��0�����q��c��a���������x�f��Ә 6��Q�5z�(���#��(ů+q&�ָ@vR�b���\�ҟ��ƌ��|�0�.Q7^�{���(2H�x��ن�H6�5�eh��Pžܨ2��n�4�ZD�98���>�ON����Ѓ�P9z)��+����C 7�N�`vq��o�a��M���O���RÑW��A�����z {%L���A�iv��5���,Z*�^�>uuN�U��iA ���*���/j������~�z�)�A����t4�.4�bb��du��6��x���k�"#�1g�8<i~<l��ѝ&~����ꫣ�z�v�n�a���cBDP��CB��;D@DZE�k@�n)���N���w׷�]k�������{�	�й��W�y� ��:M���'[�@@h��8Z��c���.ڟA�4����.D#�y�=�7-qo!lFW.���n���neh��Ț����|I�IH�y=��]Aei�1�v���r`�3GWc|y�,��j���4�70H�v*M~��
�%��8�
}j<�p��9y�U⨴�Y!���A�`�IKECC~�B\��^�*��j.hu����jD��e�҃��|!��ou��5��I�����i�y?|Q
sX��mw�� g�s����Xv���1�P���kO��R�|��9_��\FM���Ѳq�K�)�Ѽ'`kzjٗ[~�u���8�!\N��B�~����{/TOwH˂�2�BC�'0��P��Ki�$]�ͭ҃=A����\�g�{��A.ft�	����	my��6Y j��W`F�v���G��-Y0���19�W��;�wi���Ţ���g�v
|���焼����hI��鮕*��&��4ՙ�q�Ȭ��;���t�'f�38���b�&��y��B+	�L���hc
���KR��4�31[��F��ihC��2��y����I�
a l��xa�{4��  �����G��A��������' T��$���x.�LH"�2r}����=g&�~�C٭��p����D��E��-aYJ6.��n��G�K0$eپ2��@����ٿ<�����$@3�~8��zv�=�T-xc�l�_���w m	h�Ȁ�VG5�B�9g~i�� ƀ�Һ}k�,��wXety��xbhB�u��5�ʵ	�[`]K��� ��[�%�={�u~����[�%�H5���`�+ e'cW�,8�>���?Y�z�n��+>�L���6+��Q�*���R����3��7J�9ˇ��=4%;h\&ig���gY�ՋG�?��ˤW(.�m��y�#�n�!�������`+�S���K�k���"��C/����Iq�ił�p(U�H�;��wi�jL^:굈�C+UB(%b��z�!!���a�A�4ˎ�"�5��\4����PJ��������6��x��0Ⱥ k�;��%�WL@�eg�a��a����%+
�[}�j�u�qʹ&�~�+��>�A��Wd��O����������-;���}���ղS����ؿ��m0�*�4��eE���>`6�7�c��������x/�G����3�/^���s�7�!>/��th劳2�Uf�
�X�H�Ѐ���`�"�c�Y줰��?�l���.A�=���7���u�&foU��C�*
l��JQ��y��{t~zN9�#���1k�E�6V�D#�<�����?2�Ɂ� �(�Ι��m�Cޗ��XX�ڋ�2��!��+.�z���w@c)1��μ\F繰�C+$��Ze��X���𷴍��yQ���{�B���h�K�'��M.+4V�g��	yﾳ�{���^��~	!������>���u*�[�	o &"J���{�[y1J8a��Lw�O���.��Ek$cI����;Z���Ag��t#9�@��U�HZ�̕q$?k�c]#�@�i���U����K �u���7T��>Ŭ����$�|��p�31�y�v��6],�V��(�=j��!1Q��BW��5�yk�!v���j���4 A?�����أ+��������D�}��S�9q&.Boz3�6f� Cm����N�(��;��R#L>�hB�Lc9����b '�+.܄�$�`��-oq9ǳZ_W*;CT�b_��P�}�`�߻R�������yӮEլ�>�u��R(|֭Å��(+�p�u�f�����)uA�Ǻ4>�z�[a	@��h���%�GHD]�0�R��G��s�����Z4D�_�$���E��խ�VT��H~�81p�z�Ll��H5S���W:���}$�!* >�}`�����x�
�-�rV���ſ2��;$C���$���C�@5N~�CnOPe��\�{��%c��qS'!���һ��Q��3ς����S��R���t��9�
/!�xiʕ5���I ��<�B <(㎂�if^}t& Z8[����S.@��E��pn`�wl�=�E�&K��9���㒃��1�w���T�}��QS,�"8��3a�9ˠb��.Z|�,�j���
q�6����k�u���`��O�s_�g׀dY�c���;���WFuP�ly����š��C��E'�O�SVg�3ڶhB����1ЮzJX���PHwT���;Q����~y��pk,��*�3�X��6D�$L9ǧ�V3ն7�	 ։��O9�G�3�k|>�	�g_��Y�z���������l��l��X�g�	ܙ���RG�N.	��
��6pZ��Z��nm�@%�(!b	����A���4�Ī��a�¥��"�QP�[����*ۡZ"١z�x�I�A2��ϛ@(-O֛�!dgL���N �Xbv���i�vR���w�B�&�3T���e�s����*4�g���bC�b5���Ĭ��� L��2EV���ީ?���\����L��yzci�b �<�EQ �ŚE�>���xA����Q��!g�������$L���_8#	g)��T�T�aK�����#)UB�MP���@uJ�7�?�h��E�w�}"Bun��z��]S���������N�-YY�7n�p�	���A�K�C0�0&v6V(*C#����{iq�������<�j�a���S��I��RxS/�������j�I7�ي��.�L�}��%��z,�Wj�a��cv�����a*T����
C��gB� Ŋ�r���c�)�I<E�޶Y���1�^� ВN)P��� ��Ys���NB�`� 9Q$��=��\V�$}��oQ+����1�"@R��s�Q�=�D<�^e�~��;����^k��Z��;q:F�®�rl���6�P&��W�oCp�m<����Fg)���aI�� yG3D�,��8�����,�����SkR̮K�ޤ���#9ʄ���0|-�������ٖ��_h��V7���a�W	�7��K��eW�t�P��(/� �Ob��?��iB��e8�U�vK�1�sq\SIO�hS<Y��o
8�����X����fjhT�Z�(�#I�l�J>>毙�����ep�/T�4��P���,U���f�͟[C���IQi��W�.��E�FI��C�2��'�7�y�0�1�%\��ߥ�W�p��hM2Y�)e�3��
K� ��ao/Y��B��8����Hk�+�M�8=g�T�'�1ә��4��D��%�4��i�,�+�W׋5����Aخ%ڦ��&�lDZ(iu���ۅ/_����}��|��,�\Ql�-x)-0�_j�T�Eq�3\A�4>?&.TT��z ��WT����ON���k�5�>O��}^����iFJ�eξ����5��ڔ���t���;	�������&���mJf�V��� �y��\O�o?w�PG>e޸u�n�[jNh���JI~�˷U/�U�<�Z�����/J��紧�x	��*�)3���Ya%	Ơ�+�C��D/e���7Ss�Ǿ��%�ؘ䒆�����V��e�+z��0�#��gKdNw&�X�?�T���޼G0'���a��5�	��	[���BO��24�>�uP����Y�I\D�܅�^���D����>EO���s�� K���h\ϐk?��q���l��, ���H���%����z�k�ސҽeE{���8���h`=���Y�4'�	&;=ﱪ.Q��J�F��U�ZqH6%�i�6&�|�g�.�m����p�y:�D���������т�GN#k^'Z�%Ӎ�}��lJ�Mmؑ��� C�_�A�.����f��I����gw@۱��yb�����%��_"e�Ru�}M�~a#�G���CQk���戓�t���|�X�
��]�8����vXX�{�RO�(eo�*s�n��g�%�չ�[���j�=���h����itf��gژ�흅bƅ%ۤ`�� �Z���R��	B:���p�&��b���
ݷ]���g�-n�s��~��T�����Z0]t�B.��9Ĭ�Q�Qk$�S����A�#�3�zƜ1�7��tD.��b
K(}�c_��xE����#�}�.t�~�)yU &6�ૂ� -���},�'�[u�*t�6��y�_.)��f�Q+��G�◾͜��5m'�O8�%*5���,ez_�{7ǜ;��ǯ⺱|{!��D���Bo5��$�]AjsxD{�_�@�Lz~�Pm�e5���������.�I�ۨKEH�c��$V��G�:N%9��pM��JOcp%���>��s�jr�	O�~lv����X�$���	���R�3�w�To���/]Z��(gQAzPi0mT�	��F1#]��L�ֶ��>��ḻ>:�Oql��hmf�ԅ�K�\7:�20�����
���OnM������5b��ɫ�.$2�o��n�i�J��UN�Hϫ��>0؍]�g�w�h�
J�>_(�73RcB	N�;k�b97��=\��%)�jg��ɹZׇ��r�̭�$�	K5<�g��5Z�rM��CG�-222�^nV�� ��t�1��]!�H�zS��U�bkH���v��P�Ծ�\�����M�Q%W���+7Q���?�4��5��Sx���R��dF�'�HhCH��yʝ��9�M{�+��ǅe���Kg�w۵u�:�oK޼Т�a,��ybN�c���Ki>\�N7��G	���I�������w�h�ou��H��2G.�B�X�GZW��ʪ�Y0��c_]y�űdPx�F�Uդc�`â�����Ѫ[�7���e���Wþk�R�n�x�a�/$���X����V�&�[�h{�5��y�����!�:�T��*�#=l� ��#{?�w�۱��x��F��w8K���l����]}��d��x�x#�ҟg���!��P�	y$ﰃ=��v瘘\��=�[�WL���ThJ���F��$�!�s\U<;�t���M����t^[���%ݛ���_&I�nB'�E�����0�&C}�8�-+��S��Hh4�)u[�9����%�c�c*Ĩj:%��3�����k�����G�����D���m� ��`^�OfZ�$t�I���,)Ӡ������R�u&%2!�����'5�H��9k�M"Ju�Y# ���a�_&K���q��&�xI�F��}���Xm���8A!���E/dc+a1v��y}}=[�	�k��ֱ������;}���P z��6�=S#Eho�����% �S����W������<�p�e�N�,�:�*66v{ |�=���U�!)�c�)��� -N�jt�dU���ŧ������'���6�3Ϳxݛ_9�ؔ^>J�fb�xj��
�l�m)Bo��(*���z��*y�F�+Hh%��ը:\H;���}M �)��	p�3�7��ڗ�:�}�3.�G��ҮB4,f2�;Aŋ������ϴD����Y���1�\�q�>����^�"��]� 	����RL����*�,�����E0s��}�Bմ��;!��l�c�=8՗�bd3�C�?���;^�Y�\ȕ*���y�;�O��#hs作r�[ѩ�}�`^�#.��\G��T��I���/5�U��I���˿��(NCHj�$�Vc���N��dV<VL��u�fZZ�����	�?QHr��$F��7��$��.�#��1����NC�&EL��%k�D�f���%D�Y����Y�h��C��u��!����i�=��_���^�4�Q�Ҫ�[��?��#|
u�����U
`��o��
�o����ߴ)���û�u{b���Àx�
~�䃊���t�O���r��ow��(�?���&��Ƒl4a�8�:�3��(��Z�pp������e�K�P�O�ɢ���et�����R�OO!9�X�:��'�ɣ޻+XX�G�b7ONӇ���\�)�n�:��]��8��n�<��v<�����ۊ!Mԍ��=V��&@�y��.�:B�/���L�"9ʸ%����X����-l�0���s����c����kh�ƹ����$��V�T�ٳgJk^����p�TF߾�?�`�ȍz��/5����9>�w	��,�����Ս�$k?w<��G/�h��Nɘ/�J����cǨ�C���<y�=�{��^�JxfZZ!�2U�� �֖��6&HT)ڀ��->����Q,	�t]�`.8U�{Lz�4W�`�Fs�k���*]� A���������t��_c8pg���Vzo�ta�Ys:\Oz�4��5ۍ���@��˅$w!ߊ���x���A��C��\��o��L��&���m�/�tgJ��e���^�%1���'��.9sXs��=V��
u/aj�M;�E���?x���	�a"��}�~����_j�N=��{i�p)�F8�WC�e�}JKU��_��"+kz�G_8�:�Ӽ �C�0=���|�3Ւ#�����m��ep^��d�&�C���m�b(Ku�~U�y��x����4�|��:�|M��i��ق�J��V�(X�����X@�T��-��3��I�cվ}��Tj
ڹC����{~�Č�&��5>�G�Y�����a{�^����~��8�9�(0B���+�#���Kӷop�s~Ig�譢���w]d	,�H'�~���K%v�4p �w��UB�Y�HN�El�]�1���;l�?cD��q4�*ş>E��JA�
Ʈ8��o%o�:�y��	��+���50�����obl5j��T�f�}_�� ��"x���h>�ٷ�&欉�W�~���J?���X��`HEA�n�Z�0��n�+j��,F>��o5����2P��X.�=��Wm��z_t����!�+��u�1�mϞ-EL�lH�a �X��P�}M�)v��$T�"�;c!a_�Js	z7�y^������0������ˊ. zռ|��[�����n/28F���ĥdDQ�f'm^�ߜ�4���֬,���6�Ti�Q�5��,��Q�����'��)#���i���v������z���#����g�h-�>�un�.x�����U"זf
�BHv��$���;r�����@ g��* @��)�0���7�?�0RM�N��n0	���). �!�[�|� ����>'��{ׄ\.�<��]TUCC��Ȩ����bɉ?��/"{),�!��кM��� ��BYY1����;�/���(�\胧��ޑ9lBq����Sz��e�-��P{���S2EM1}�v�%��wx�g���t����ȱJ��r1gK�E��:�X�����~-*����-Mڲ�?�ӈ���-�1�Qc��'ҫ&�e�:V�
('\������Uh�SSS�"""�O���Pn��}0����pr"䪵4%Ө5�$Y������6��T��/��H��� GQ:@ Z��b��K-��`8z�x4����kاjfJQwg�DXX���-q��)��e��g�aZB��:V�O��]��\�p��n	��������ƶ����P>1�����Ȏ�~S�b�ݧq���J�g�O.9h%��?�{m-W�A7���a�r��$\lc,�$:�tH���y��=T�F��b&�+}Q@��p�6_5B��?��*<�Pf���Ӏ�@Eﾍ�o(1��,X���Ƚ��~�U�r��cP]ՙE��b��;k\�0	��R ��nX��W�^8P��K�6��FO�W0:�m�
�(��S�y�ĉ9"��s.�C�ڪ��j����1��W�2p�m���� i;ͼ;yPn�Y��$畼")T_g��r:~dD�q�U5�9�~�����kb���p���3��I��p�Kw�'�@F��:���n���0�P(ˆ)P(g��a�̂���]4l��Ch&�/��Mem%GG��`yj`O��)� \U	hX�!J>
%|��.��f��[$����������*cdd���� ��9�%��<ŉ���]M���"���U�4�u�=�&���������+����!�g�9��̝�2q�V�;ŝ�(�i&��zHT"`��7�a�
.0�W��bW���U�
Ǚ{Ec5)rh����m��S1l�C�y(7�	F��DFd|��'^�]�5�XQ���Cmi
��1�HA�ڼ���u�70�Vo?�!$ �?�.�\��ʐ��c��?�ˡr��3����-�($z���;�nb��k�Y����u`kEkρ���V!9{�{�?��-�xЊ�ohs ���4�9��Y{/�^�C�h�Hz�L�<��29�=����`��*`��X>¡�v���J�����2�`�`rK=���>j���M,KKFHG�|D����4Ӡ\π��O&��"Go�,GѸ|���N5@R�,1@KAj:%G����}$����6�GM�0)@���Mi��*����L o��7 ��|�g��!���w�V�ϳh� �k�/�h��yu�/�y1%�+��U�%����y�!Ss2���;!$m)�����/-�������������4Y�Y�Yn� ;Z6����V�8獖�9[& ����E�&!�����d\���U8a��е���ۗ�k�Ǘ_[��2�{��9�k{B̓�+�m�4�fxc��uT�y�'w�T�3������R|��'[�6Q��l�ۋۻ
��#�l���la���Q{��J8��GC����,Kͽ�����5��� ��p���B'Rz���5��	m���VKv�̂<Ov�٪�M��v=�T�P8�al
%��F��.37PĽhܰ���z��2�Q�;�+�[E�ccqXY����|kʹ?P�Y��� m�y�x)k��2�P�޻�:ş�R��`	'm"��<�����>�!��AXg,K G���b&�&�%w��>�Z�5�X%�d�ܪYgSJCD�LdP<p<=�����x���VZBv�Xv������lᓈ�Η��R����&�����{ө��[?��'���,@׬�!Q&��tZK��L�R�i˘"G��θV�0R�u�{a(z�#�,�%��Bl2rr4�s����=&-њ�cMt`M���`�(f:rđÿn�Q��wH�Z����a�3r�mY����	x� �*D�_�A�9��M��	����VO�]
j�<� ��g�(����'�\?J3M�BѨ�?KK]Ny��=�_p�-�z�)��`:�)5��ʊ�M���Ty;��58V�����n2�Y�V�����p ��-C6�)��2��3Gm��<7�Q��<��Q�d5� %��UIQ��
<����r��}�B�b�+��_��I����q���9��>As���g���I�%�r����ʂ�>PK
tHj�e�f�
,|��#F�zb�<�Maǌ�X���+��)�3�_�~�Sq7Dh!#ƴ#��_��#]PS�^sC�`�m[G��1<�ӽFg{ʾ���'�
�b���'b�^a=)�6�H�ˣ	�C��)�I}��y�n��9��cpCz:|�d��"zml�� c�X�D�$8�s��*f��k���~����
�j�����O�&t��8w!r���ڡ�u�7
/�c���h�`)�
��WԼRK�<ovC��a��G�"�S}$Ih�מ$H�h�<�?W(�cw�\��;f0�n��Q�Z)��W;Z�J��hp[w@bWq��B�EkY�C��
��X�o��7��h�cg��.<�|)pO���,�6bAduƙ�]I�����i݈>ev�>��s1$�1XB�!��'�/�;�-`��>��L�o�';�+d9�NqV尫�h�����LU��]~]����4D���$-|�L���t�|o�yV�"̾^�7z�ѓ��c�g�ѕ�N?3U�W�]���m�g���D�mbw�˃����O%��B@��m#�[$�zCR5WM���_�,(ދ�{nmv�r��$��i��?w�n �]_d��D�>u�՞������6D�����Ap�!�[�Y{3��,�|2��JR�L��=�ި��EX���,�K0h���q��!��ZE��n@;f�/V��C�b;}53t�Sz�l���)t���0������35�<߈������w��,6���O�&*Ϳ�\TS(�Q���Tr�i+CP~ŭPn0�݉1���,8�{�ը%q�}�1C��p�E�
|=�5��?�j�0?�v�mҋ�6�#��b�X�0ګT��$4�D�Я�@�������tGɇ5�I^ne��祈O��H�+����b*���ma���ZmZ�*�F[�}ۚ����蝆���7�J@+֋������O����k�/<�LT`��c�6g�﹍Y�����`�R>�cB���׃$�F�{a�3!W� �p�s��d�]����ⵐ8�Њ+6�>z�ꙧe36���L¢�0�%��>��Xu�:�=�g���єG���P�5�]]3'�C�K�Y��� ���0�;Βf�*b��E����<����.;]��Ir��n��0�&�g�D��y�eX�{� e,q���[�3u��ux͒ǌַP�7�p4bhQ�� �E�N�����l��R▋�t=��D�=�ZLV������ �es�HD
	��F����O�Ҏ��C��0�F���Tb����e* �"[��5j���2�<ѐ��y)U���?�������D�%�R�A�z�Uf��<"犿?cmQ�e	����d5F�!�h���w �!�ˏE��G|����k���`�&��ί��/`�9�u���m;.�V�m�����Iy�A(��1��y�#R�O�d~�C�%����A�I~��2���9�d��'�Ѳ�]���+o��������`��D�OL����X���ܿvRȩ�d�6� �n4��2�ų����#S~�J���εb��v r�tu.�{��O� �A4��r iF�o�X}&�:u˯$��n�^���'s�w&���S�Xz,�4�� <=��x�	�!�M��Xw�;|��^��u��2��:�A(�Ä����c
�z�T���*�8�t�Gqc�
��� �@�H�!���x�Fȶu�u��Yr.�е����P%�����:� ��Ѕ�#��N�X+��s^�}.A�%I뫄6�r�C8�[V��xi��N���CQv
>|��>���Jbu4�ֹ���ua<��-₽#p�X|!V6���ބћ��`��1�	7��kɀ�|��g�dyc$M�N[��p�����%-���g-p�z{�C��7���K��%���Bk������Rs���Qc'$�I��IXAF~�{�K�g�L�G�V��8ş5b�9�O�3װS���np�L�q�q�4�B�\@G���k��s/��$�m����}1�b������/a+c�.��hT��=V��M��v���)6�����y��%��8.W\��0�\/�k�7� g)��������I��X*��8��!)��[�o���|t)V�-���O��#�w�������*�*|z�C��Q�ķ:�̧�#����W�@�Ś3��2~i��X�}�������i׏'22\`�ۑ@��itQ/)Q(�Ug������oa@�/ U[{�yM�\��-����2��i
�e͙x��K"�g�7�7+E
����'o�v�����|��w����Ӻ&��z�	�	~k��KK�&����w�J'�}���d�¤h)L�)� ?L������&��� b���k��wP	$���t[߯SM�7p���{� JA��a���\\!gn�Kј�uǪ�{�N�!�V+��G��~h�����f��THq;�B���s4d�2�����@ȋ�¼�`ȇ���.���_���x������`�%�\�z�lm����8�F ��|����TY���4�  ��q%�F��������u��D�"�s�c�F�~R�_[-���3&Yu��0V��8h&��+%b?�^����� z̪��ֿ�7mnA��7]$r�8$*uD� �E��BCm����1g�zd8 ��ܛ=³D,�
-���qH��N��;�߲8Ce\���/�o�t�Ӂ������{g1Hh��sg�3�
܅ѓB�D֒�b������j
4��ϱ���_2�Z���
��\l|����7�ͼ������}6��)�x�/�+6���=��aS������w�WF�S��,#���6���g)M�n���X-�|��|-i�0(��y��Hј�ÄNq��ؠ�9�/s�g�rQ)��&�-(4�, Z"kjk1���*4G7����(�w٘�#��1���V�&��m�!��]�G�)
�Y �5�lG�_m59+�b�Կ�1��J��v�;F� C�@��݂��[y��%q����R~�g�A��1�"���������k-Cq�1�ے���x�jn|����<\��F�U�}�Cvv�L,�80>��k��iA��'Z��ۖ��N��ߡ�9��3^��f��֦�A��ޙ��I��&��	������"�YE$�_��?*�$��a�:	�Ǒ���T�k�:/��hM�<�����6Q^AxCμ��� O�R#�$¢�7{?g_d+�|�*x� ջ٭�5�8%Q2T�>��2�BD��H쟯h�N��]ɣn�6�/�G.���[� �a�5i�j~޴�K�tO��M�r�䍷5��X�J	��ζ������ ���)�#IE1���7�ub�#ڑ���Q]P�q[Cn�nJ��W��U�~L�)�� �8n�WoA(�U�&Y�R��N���"$Wd,`܆�޲ۑt4��(k��V80&�Hr��bޡ=��C^�'��g����nh��=�I�w-��W����N���Lz$�[i��lBq���VI�(/�a-���]a�!/51я�������鋎![�;���q6u:�uJ������jG�j|m��-#]���'S����g�*�y��H�{p r�����<��f�����%�N�áU�=D\������[k쪝l��O}#��&\
�G��Z��Q������� ���q��[��H���U���!��ۇ�����m����oÙvBD�%��{�cK;�����ɇ�bM��t�`0�$�r��?vǙI��!oNV3h!ȓoUJ�������A�A�HXVu���y].&F�I� �ڂ����
X��,�D��e�<���[ħ���0�ҟ�s��s�o��;E5\w�8f�[�~� q�ְ1Z[S����Jπ�:%�����ʃcŖ�=��y�#$���'�R��y�� 0��g ؎�\A�m�'� !MN�����0k���@��~�j̒�����.~u��,
Z�-� ����5?м���կ��?v?��3�����.q[�~)u��|�R��թ:NI@�@R�#��I�Qqܹ�4�;���"2�e�h����q���D��H��K%�]��-�r�������� 3��W��3qU���s���ℎ�?М��W�R�~r	d�-�����}c����}��Th��G�1N�~:��v��jz�D�&MC؎��Nz�)���HԸ�x<�JpV]qFN�q���)oz��h�S��G��+
_�+L�w�W����o�#$F�wr?s�O�B�/B�c"�x�;b�������D�ep��r�1D��qC?�����{U���͑o�f��3^:Q��>�u����>�F��&Y��鿁8���8C7�DC�xMD �3O���P��� 7-��mխ2_��0}C����*tt�6�����~��~>��t+c�y@+�̋V�/X�~ո�(b�*O�9������}��}�|0�@ӹ�E������c�3꠯L&L�v:����g'=�#�R�S�{�j�l	��¢������F(�]Y��� ����tG|H�����{ ��Oe�;% �=I'��"��&F�nD��'O��행��w�Ç�v���~�ӏ�e�GHy�%���eHB���+s~r�3��q��(������8��(��ض�>`�(��,�so�&m�9�}�X���.���ن޳���/�!��62�������"�\he�>��`TO����$���H�}�Xy�;���}р�M������u��'���ۼUE-7�\~O|�W�����n2���a��Ȗ��ne��=�^-j��m�����
R������\��qT���#W]m-����"���$%3���a�i-'ϻ�c�9���k���'��b�����5���|�� $������P��⁝���6Q�����c���W Q;}s�-C'��]��(!�E�o����;����o!!��*.�h�0Ƌ/��Y�*����}�g�6-8�V���6wb��5�0���ʎ�`fƤ��P�+��  ��h�ii�^o����%����7�jlw�@��~U���;(�?G^�5-{B���	6X�P�;H�l96�E�y�u�����1����4�)�0^_V&# �.b?wt,]n�[{�Q~�?�e�N`��U����A�ցL/�����ڃۿ�D��-Gk��ޅ�x�3ݔ��ֱPv��^XR�����<�b��n7�!��3 �B�*�{l��GtU��)�0�(G��n����L��o�/3E�{�'O��ovX�tK�� 1.5��dJ@������|3�Q�e��'����$�����������р'��������w�צ��?|���|Z_��~R�H%Y��p�׫/���%~Z�g�j���O\9#���"����e��0~����=�a6 ⤧G���>�p��i=]a��҄PhȆ�I]��;���N8��;�Ib��*Ե����w*>j))�����[�b���rnw�|ƭ��|f	�9���<���]�i���}�:'^�k���ӂ���t=����[�6�5:<ܓ�jer:�e�Ǐ$���6P{����ڣ�s_\�G@�V7�]{]�KIM� Ӿ�y�־�ѰO�c�)��ԙ6��з5#��+�\_F�BE����p���-�|�ҷ���[Gǟ��-i�=UlHNNN��m�F���uB�/�mq�Z�|�P��U/g���p>}��k��bo��|sWܼk��a�u�j�[0y�Jb�٨��C�ps�l� s�F�sA����G�`���߈��h�N�����9�<d�+X��̏`�㇤��{��p�I�o�f�.}��땛l6;�E] �Ì���X�������
���hXkWXWF�^ ��%�w�r��SeO����L���C"�xkN@���)�@\fR�_{|�p�%���s�>5�g��:H���2/ȓ���C��㟠��x߽̓M5�Ҥ<�g�{��e�f����m+����6j��?~]������� �c�ڬ�_��L��g�ϾFa)�'﷐/�V ��@�,����s�֜�?�i$�ٝ���P�_Y+L��o~�V���;��U��b.ݍ =6�"��h�̅�5?�?Jf��w1���TM�sp�P��3���+��i���F$#`+=���%�b�(��|��m���1dX��>S�%����&&"J�*�vb�&��ue��'�>���%�W�NDDt%F���bӒ6r\9+���$'��ÞUu�]�7��ůtyi��K�w�?(�@��"� �P+���<=��z��[TTUU�?=�S�5[��!Q}�(�!6�s�e���>)���jw,ׂ~���B��?��P�5��0�
�
���y��?:�׃����˸�{�c��@]�Q��ű@zm~=�jo��sW�Q�E�����Z���!�}���i�o*��6���ORs1ρ4�pE���ĕK=mQߏ~:`p��fz?e|��O�W�'�.�*�T�_sb���2�)�.&���>����N��C�*
H���$`Pi�����N��Y��,���7\�DXNp�d���w�gc?��a�,//�����P��O�wD�qT�G�q���4p�~Xۼ��hܺ`_P0[�Kw]�ة`9�k��@~*.����4���}O8�����͓�95�&���x�j����ն��{�o^�����'9�>��
��(~*�W'�T�f/M(����AwA�/_����ӓ��7_������k@����/-��UU��M��̓ *�k��m��%5Z�O��ڝU}�D�r��W���
� I���{�{h$=ו�\���2pj��tߴzكJ\��u ~=��ICe��a��Ύ~�l��|�'=c���S!(�9E�S��(0(�~��NQfTK���i�V㬳��6���˥Tr����-	�P�n�M�G�{(��W1��Z�n]�t��ɿ���� a�o-�K����ⱒ����L��B��"���˜7LC�K+p��������'i�ΕW��u,�e��t�����`��Vf�H:�ť�y�����u��䚟�L��4-�����4"v�;ؑ�Ġ�WMy~2���4�}�%�?�� b.����s�.��?�E����M1���������	a�k>���m1�k���!b����E�_gIMȄ�+�f7^�waX �} �g����: �hk�t����]R"( �!�%��)��tww �������{��Ο:��9{���߳�F!IM��c���F�L	W�U{�R��mn*����/�VxJ����o O��V�������G�����.+�߼����Y٨9���L����Ń'�U���	���54@��g���6����g���Oi!Cc����`�=�`��:�ۿEA�6]n13���GŎ�������P�V�@Ʀ��E��0��/�"pR܎��$�c�eY�#� T��O�e�*�(����y��#C9�uy{SE^bW�)�M=�?��F}Q=)F55Q��ھ�A��p�T�o�3Sl��������0�g�z�5�6o����(�?�d;'i��ׅ��?�!�ά��d���:��x��aWw���A��J��/I���l��=KI���+8mS$��6���� 5x�B�V�ށ�ΰE%���o�"7k���f�:X�OJJ��+0~�ջ���������V6����Gqi~:[[��̍����m� ?��{m	�<t@��f���ԴT�8��7B���K�G�"�#8	�ߍfn|�7�����P[����PvJJ��98�(B.X��B '()a�ei��u��<�o��\�<�����i3{
^>��mU�щ�E�0e��\�	�p�~����*���r�_$҄��i�������E|
{7�4�p��v��@"ѻ��%7���(���v�@�X�����VX�X(�T��� IH[����4�+2ݺn,m�繕�z��ϓ.�����^���#A[Lj��Ŭw��rr��R���.//?�e�RCBw4�;��&44���*@����������K�������8j��������,Q�aa��Et��7H�ɯǗx����|��il��_!M7�I� T�>,��'dC.�
�����N�0$+�C��Ť�P�=��3����.�=&��v zp���"�l/"��}�Ru00��P�iBgR��֞ިy���F�-���z{{髕����@ԯ�f��!z�簭���_� �+��0~l<'��_@|A���S��k�7z���:"4�E�g���)�kWkqq��Y�P�]\!�_�FHY��_6�4� PQ�nηoݛ����\pZ���	0^r6M�΋K�\�g~���@�ʩ�A�sd����P��ξ�c�355ͫ������|NW���w��@D�(뮧�+5K虙�s�$~M�}Gy	Z[��܏����B���yUU�
�៦?;56��i��p��#Ɛ�ll�OHJZ��g���jf��Į:7�s���!q�
�h�*Y�j�=#�:L(�oMk}�	�]�jk�ܟ1�.N-D-Hʦ�I+�7|�5G��7����zOv�ף��_�������'���95�֝��K�K����/<5���{�H����Vu���U;~a:PD���Kyہzy�G��������%%SN@$�@"Rq��]���W�8/��Ƀ�bҖ^[��@�Sm(3�L�<���笯v ղrA脙C4�k��V�֓ �j��˟ج�(>pns31��N/����wL�'L"����ha�uݹ�e9@0i&5�!�C����M�#����巸�8��P�Ģ�Q���G�@��jٴ�|p C$��%��Nj�C!hI.�%�=Dg_�ƒ�*���)�^�T����?`�ʝ�6N��y���mX�=�2.K^��$�|8=�!��Ƙ4zU2���]��g�,�JD-��U�r������6|4z����F����E���Y\WY���P���+��a��d9x�����7�[�z����]~����Y��ȗ	��?����#�?���3�V�_�^���8��8� �?k��*z����sw��j�s�;|�T�᱒/� HZq�x�r�}��"�C�����Ra.�*��]̒���F'&Pr���D�ϟ?�;�A�:�;���G��CY׫'�;�OR�1�-˚�.���n��F�}�#7�<�wc���g���WYY���)04>�L��o��w��5�|�
Tt�b=���<��R��}_!���Bݾf��K�78��O�H�������:kky��*�ę变M�0EΐZ�/��/��A3>D�y�����%!�t�D,��/ ]P�?6x�+ $��S���>j�k;��E腅��=��c��"�wܫ(�DH,�D���䰘�-����;����ߎ0~	��~W����3/��-�d(N@��CNE�"�����i��w֩���,a=ᧀ��4�����3�U/`o�0��Wv�de=�l��LX��C8��b�=�zB�g�^�����π6�)�ӅUc6��EU�ր � ������5%����o��-5�������gL��{J���t��d�KU\`�Ͽ�;��:o^��Z��%��\�@�.���D6���vHW0ƾ�X])M-$��&'?�V!��^7cW644�s��6�u�o�����K��1/��	�G����a�);D�b��������[#���F�h��3q����b��񄅲�+�E�c!�(�e�k��;���|�0��´4�/�_��E�������[v���h%��wv�"�����e-�;��B�<$~�ht�rk�ю4�R^��|#�Ԉ��{�c-,��E&�t�4k�>}���Jah}
DFtFR�c&iv�[���8E��Uw8[s�b���{cww~֖����Pg�xJCEHT����[��7��#��{���zǦ~)���t4hΪ(BN��}����E��|��\7E�i�gA� ̙E���AԊ~����r��5���s9���A�'����N
�c\jj(���mn��XY11��C�F��i37���7��

���5�@��9�/,*��Z$�~	���T/S��Y�:\��n>�#�`
���'�������&7.�K�`�	o��TZ�V&�����O�ʱ��s���*yjUk+)�RF��x	�pH���$k��j�3��6�I]}cK��56���Es �&L�E���ambF��P�c�q�`/�ɼn(�m�c��i�t^���j. �~�B�<<<t}z~�\�/@�-���(�.Ǻ\�)������I�%:F�ٻg�ǵ:8 ���[��rh`21�\@���J$`�����	~�F�����Mݜ���
�ǚ{��k=Nl�44�{����'rG��掵�)�a6�}ۓ��
 �)x��C���J�6w0&Y�Ȳ;�j��Ԣ�W ��7��yu���Uxu�\�?q`�������\��P�#�����2���k)��N�:���G���Ym}+Y��u�.����؝pZ��L�L�V�']d��Z6��S"�w�����S���9q���w����Dw��$�s�jF���VU���\��������J!�����(��͵��a��E�}�������"z���`��Q�;U�w�cL�f>��*��q��Z������WLg���n-�:P*��I��D���7���t�f�<�~46L>�ûn���,xz�1[��΁��e���V1�'#T�	�[[�f���q2��p?wN�y�@�3�uX�Ff��b�:\VL�1L`H����=0 �+@�QB�������i�u+�TG������A�#I##XP��|�(�п�w�uCh ���K���g�d��-��OS��2�h�䈮�a���B\ݨ�B���
�bYH�x�	�O?Y�[�gH�iG$��-�9Ł�# ��""z��B��
�M�Z#|��{��#�K0�hh��w��pj��չ���@A��p' ��˸�� } Ox�7e4�8!H[�UX�ڊx<��o��~�F�;:#iw֒P�1���R�IJ_�T7g��p
0HÒ���OԳ�	��|=�t46��J��p*�̵u����4�Hi��Æb�Pӿ�4�]����K�45;�N���D��Y։�3��|sPDݫ��F���\��5$S��G�dNRCYqD��w5D>�I�Z��F�Jf�*=ә-��wp���:������S�D��<�����nB3Du<fAYe��ܺn���f��d� �w���no�|�����|�̰�Ut\6������꣓��9:�)A�\SSc0��Ta<�k��F�����n�/
4s�pA 
�]CP>�*Dy ������Osۣʕ������YB�ma`LeUUl�`��Ga<*L;�{D��Oc�A�w�-�."�_̥�8:;��x?�ܜ��n��/X�'�"1��|��Z�)˓*~�v 8��?�xN����
Ox���T��S=��:3�WG,����u�FM�Y��-�����ù��Ox��c��pp�!m �ZwwB�z*Sf9�bl�E��qI�z��Q'	�� �3͢p?��rw(v,P�*+��`�)�G'-��Q�k{�LQ��S#�>]չ/]�7���ɖ�4�HŅ���O�L6.`�直��}�0��+v�#m�Lk^�M3-|�$�k����%��lf2Je>	�⢢.�h�=�����ނlﰃ����	�b�_�0^@
F����O�#dGv%�̛~�GO�Φ��N-��jl�� �h�y~n����������)�6U�iz�z�٣������ݫ�l��9�1>�&S��àQ�/����^
qQ��hN
�^-1MP0nD�|�bC�{ur��ۓ���	����7aΰ4�~��v-��{� ���|���9!��H�|w@+V����K�p�
r�����FҸ�B١l�&�v�x�ُ�	j��sɿn=�2�m���i��N��e�+TB?;8^�����!(�j���D��Tn�;fd��0[��@t�R���9?����b5���5�҇�-5�\�����6�9!NHL�M&@}������Ҧ�i�JX�h�;��:�c� %���Ǌ'����f�R�d+����S)�F�u�K�|z<.T��k�+�v�W�(�?���-����|'7�t�c��� �a�pY�m`^K������<�.W�ǝ�w��aI�}H֮��H"���:�e��f�f��� ,��"����6����q$��9���v�[���?|�fQ��Y����E��x_��wY��Z�BVnk:ܯjy����j0^C�8���0���pX����,4��K�?��t���e|�ma�$�ǋ��O�$�K��z	J�:���-�X9�K�ds���$b�;22R��*��X@Xs!�j�O�2@�3 �� �R���'B�w47s:.�>k�7��tM۠��6@e��bbcs�����u:�adb��{�)��#hT4]�р��TEb�Vһ=����sNS�����W�Q��C�)d�p�y3�像aL��yї���}٢���6f@>�w���IJʿKD� �؍����I�@�h<�e�C��Bw�2|>�j��o�Ia��^QQQ���!���ʛ�W���r�e�|���c���"D��D�������W#fq�v8:y%�I��XAI�,�ko����ʼ�6*�� ���V ��C�虦�}�.�?"���w��?҆������M��6��'j���S0~g$��t��m�!#��N8g�N{o_�-�qN\y�L[|���@��/q�W���n*�<rq1�kr~ޛŰW��Sƀ���MMO7i�y-Ө�5S�ׅRz�=�h ��g�1�Xfi2>��U'�~�]�eKg͘�ԑV����o�I�q���0ΈKH�o#6]LV��`5:2���X��j˗M���v0��}IDn�|��B-���Ilm\�1��?D��v�u��M�����p���������ln�aj�kd���Eag�P��2wo�S:�\��3ׯ.��?R'�y�]��C�����h"f_��d��c�j((�h4�Ӭ��
֭�P���.�	�:ˡڑ�o�NN����u��r�[/M�W�-�.e�4���'6|���e���7��.˾T!�Մ�����I�d�&�����(�Q�j׮);��V����{� �o�r�ɔaŏ�Fµ�5�V�%�O��4T�_T��E��{�lnv��p��ҿ�=oC�F���&���Nu�(�7܆*�EoXN��7t��\U[�9����O�^���>�lWp�F������B��8�2&E2{e�č�ݽQhZ ��`�Db��,�������-��P�	���d@e����Z'|��i�r����13.��̂���j_��*�0����.AD�l������nD��r�If��w�jR||�d4X�;��~��8�;;�i�[�)aVx���(&t���#=c����M��AK�a�2��1n��-:� ���6����H�y������>��V���O�|H]����C�]�r��g<}��%�7���!%�R�ǁ�Y6#A�"�a�D:S��̂�+<���/[��F��8�N(4+��п4��,3Q��c�_v�F�;T7cQ�����_�{�!��+�ʄ����j�1E����V]pP������'�<d�@�����ؓƕ�@T����;$�l2�d�7VWWO`���32$ݥ�+R��T��X$�9ꖙ�ˬ2z�1Yl�߽{�g/��*Hz�.��O��L��xDTV�n��!9V�)w���JI�Ϋ���8,F����"�ܔ�뽑D�u.l%;�~�,�DDR��-0���O��Յ.�Q�|�h!�K��I�����y���%Y̑��T���5��5�O��O(XXR��X�����VW�}\��~*�0﫶G�� ��0���<��a�ɈCS����FmQ�(�G19�^JwO�kK @���ttvĲ6���k��`Q�%}f��||�0�?�dUt4���y�Ɵ)GCh_*���u]cOR4��İ��񂙓[ϐnJ.7v�IH��(|��I}f[7n&��=!!aw����-� �/&��n�i�.�]d"ڮ[��U5e
�u#'$&q��~����p\g7uu�=CE��߫�����P%�H��א��R7!��ѱa����rnAA�R�����r��*j]֕�%����ѦL߭� ����i#�R��'�
r;��nA������+�D���s�}xdǑM4��ęE;��.mX�
��ε��\b��ҏOE�$8�%rf�)��r���5�x�?�|��I1�����fF���󃉈�̭K΀۷�}9mi�,�h��d�)���Z��ɇM�1e��N'��*iQ�-u����5nθ���L�o�sӫK��\'�����`�5-�%-�G5�Hi���K�����91�����|Y6�j��pbX/X� =�~^�n>YG�x?�g-���<���EM����+kE`꧷��/v'���q�!�-D?����X̑>��v=t���0rʢg�.�<Y�) (p��C����?!͊ML�!�����.��Lj�'A7�������5:��	'�̈-@я��������|��%'k��Y(r(4�8������g'7+�#�{������s�8��߾�17X�	�Z�i�,ۿT�J�~uᄺ+�� ^l?�����A ���0��E�S�ez�G���������L�މ�,
R�ə���+G���%Ǆ���+�����%XƧG~�&A��Ϛ�A		8����7' T�r�1�p����yejj�rQ$$�G�F�X�"n��$���#��
���Y�:e���+�f�Q~6���L�ug��`�?8D<V���M��e��!�6�"��%��!;�o^������r�+��}h�kN��B�?
%�nJ���Ad�����9�������BZ��>����	��s!�����t_6�=�*��S{�sY^^��?���ޞ�jW~E>;;��&����]�mra�����R�����Oв�T�y����66dGe�z��h�ֲv̢i��^�j�����x���?B�����<�.a�nF�El}�v��l' @��xs�j��h"�WD��5���u+��1E��Y�3�Rm�������|6��gJ��S~r��܂���~e ���?l:��.⡹�tٮ�`bcbf����JiLL@����`�]6"��rC�F���G�v;ww~;��ܪ<l��a��(��s^#���2�ʪ*��~�B�k��@�c�w��l/�[{8jx�=ҽ�q�k�v
�����䶖b�1�#����ru@0>e�õ[��*��v�p��%P����o�H��|�����lӚ�����Y;���
����;�.�w:��T&�����b��� 3.���&UkmOO.�%u�{�e
�F}�
��i������;��yN�.�˴�\�K�R3�b�Ǻ �)�ؾ��� wb����"Ep��~K)P<�W�k^&���օs/�N�3o�R��R��T�WJ
�d���>9

���:ͅ���6
Pf�T����6W���m���5�+o7� �fI����G�
�3��wt���VoV�<b����,�.�*��#��o��y�
/:����4���c	���b��~�=���UR��@5�B��5::F?6����}0�D�Rk}dT6j�w��׽��<�)��?a��*���Af�K߁x���?��T����G�90m�/,TWW}���\U���R���;B���������Ōxm8$�
�8�Hl�ʌr�P�G��K�)�����\�nD@9}]�P(��X�K،�����&5mi&���#f_�,��i|�`�]�n�$>�E9*�&�P���A�`�4
i�Wt���(�V��	@�/sh���\V�����T�@sD��ml\�3tՈ��6��yA
V8�e	��O�	�8UΣ�}f�>��<<���N��ޅ�WXFE�I=}58���<�9� ���yrbˬ�A�g�6_GM'�߇ |��Hcg].`��Fδ��-W�t�#�*�X!�N���ff�jm:����B|��G�| "�Ѵ�G�{N/�Ό��(V�z���&VVh(n] ��]�އr^��vg�#�
�(D"3[8!̬ y�����O�w�-%����`�����H � ��G6�z�:&G�����C��]��v:E��~h𣖖@Q6�d�ŕX0b�F����ffcF���
<ՙ�A�K�O�^� �g5ِ|�'"�JKKSVSqO }�����c�EMc��򁊲����eu��Zg���8!`V[�ھG�ܹN�8(�x�pF��'�H���^
��{�W˩Ț9����ssr(�j"_�JIr�
gc��F���FSۻǿP��HA��5�e�c��룦*~�|,�� ��Ќ9$44IK�"��)�k���2���%*hr�_l��0�]_��*�S����n�m敕�u��^�,.�،���?����JXJ�q�V�	њ�ߒ�RcIi��o6ӾTlrZ�_ƿ�0M1��	��WtR�z�����In[8��Pm��<��.��&2�P�����c�՘����~P@��.sc'tDQ� Q��a��gl$R�ѕ<O�����֬_�~]��d�h=�v"lbdܞ|@�G�)W�L�jy[HP�|�����ZϴT���h�P��v�Pb��˘�r�9��f���c�DL��i;Ȗ=��ֳդMhu=w��W���`&h���.U�o����pd�"ka_�2#S4��:������Q�r�#���/><o��h��v���.x��p�y��ef�܌�u�z?9FV-�-:�W����tBv~��f4�Kw��z��1{48�'�ˊ��/�,"ǐ� �3v`�g��'l0k��O>���"��"�@[y3y�^�[�Z폥r�/y����M�a�a�}e�O		�:�̆W���d�݄�M�;��Ґ�GI�.w��� �`�(��ro���,.K�vl_��;�u�_fu�E�?��%'���B�.u�n�z��;`� �G���Z������p*'䚫��V�=0��&3#�oa+agl�rM�YI1ٚo(%�Y��F���koe�Ʀ�������;��-`㡻��1�a��mл	je�b_���k��	�}���L7��Y���QS3���
4j�T���w�lTE��D�Yzݗ'�U�X� &�Xkl�zl
���Q���wD2�i��B�JJ`´fЍ�n�KA~xH���(�	���1�{�����<���&
_7�K��Ʋ�p��;��A���_���n�a�ɜ/AP����Ϙ�a$�!V��X���� 2�+�1"�!5����97�N)�Y��JQ���;m`����B�k��F6����Σ	������Hz�f��q˵��Ӯ1l��<d1H5����.Z?%2���8����u}�W�
�2>@Qv\嗦<���8=Y�g�PMx��.�s��R&j {	Oz>�g�� ��?Z�����p�<��D>������9X)�*�����`N�[�>�\GS�������Ŵ�M_���wFǆ��/��R/j}Ȓ'��Ȯ���SЗ�V������z������j������ζJ�)\�hx��F�#��А-�D�������4h �U���0��,qݏ�q��g��lT󃧡�����#zt������z���嬪}�����$���h��
���g�'������l�g�8BiQ:�E"�!�4(@��PƝv^v�ʿ�a1�$���/�Pv������tU�� T���v��)��<��+��XΞ�Y�.+s�����Q�����u3' ���t����S��:f\���
��
66�R�6&�#�V�g�]�}8�d�'2�Lv��2+|���!0ɜ�����q_C6��:����j����څ¼~��;p 	��F����ܜR���=�!��Pc���.�W��t}%�g��|�����G	.J�^��_D� j5�=>�a���RzϨ��#�=�H���ޓ�}XYy�B�i�-�{����z�:ĒQ(�dREP�rG1_�� 	��H	���j��{��"8&-),300"7;*
�g��t��邬�
;�_
�l�q}||�'>l�_{gkp
	E�`w(�!c`UˆuS-ϙ�K��Tɳ�ٲ���ѳ~d'ܼ���k�6eo؟6�s��K'$:=;J6ͼX�79�/�l��Jii���E�>_f���	{���X���#S�jy��]�=�܀�TfHL�?�p@� ����}�{���A��W��P�6+���x�������`���En�b��<dGg�	����ږ���=`M}����̲����c����`/�Y�%.!��RT�F������8i1�i��
��@.ET(�����c���p�;�$���8��uJ��Q	��)5�����8Ɣ\�8#�����!o��u>~���599a�)�������6<��AB-��m���c�R
b�nt0�ٮ���<��~&���� ͱ��cc��>�������Ϭ�[R"o�u�u�Qgg�r>�V���^�3Â0���n�<<>>~w *^��u�x���+��%�,�8�tt����D��N���كdя������+�ppa�<Ŷ�GԌtab,����MJ�Ŵ�h�ˬ�
���RU���-:=��#�Д'
J�j��G�Y�@�l�u��L�l@~���&�@�����ܿ�������K��2v�N�h*��}�J�P���c� �M3q )&-�o>>h	퐉�XG/��e`�-,-bSB���S)�o��ͬ��$�H����Βg�6���B�3X��Yvݞ�)@�Ǚ^���&#��2}�C��brfAb�D���M�ӊ
��3K�,�ɯo�4�i��x�=!ƞ2V����~��G�z�Ѷ����Y�
T��9�!�+fG~��/��n=ao4Z�����3^c�"��^�������YXZf:�����JJJ��Åc����Hd��]�Y�Sqb���a8@m�\�	?4P��ӊ6o���#0�f�|��H�I�;��z��&����F/:qY��$���-�;<_L��l��55��_ݕ�C!����p���t	��t�T&���� �xh�gw� ��U�����V{���e�]ޔE��qK���׌�|�i���''lG8��YCt4f\\��ׯ�z���Y�~x|�����O}����8Yn:��zm~U���W&�ɻ�����$�B
`s�B�aŏ�|?�3Z�o�\J��6� P�鼩O_���6M9W��V����<;?X�0�<��I�f���+��^��x1���K+q�c$l���ι�S��L�¤i�uk�b@�TV���ye8��Z@�<�.̳}��>bB\TLY�nd3KX؏������QI6�N�j�$>�)����v���B0Y��2bbIKy�nCܳ�3CCC@�Q"��е�b�u��W�~��(J��R%ZFŅ{� `�?���R��X�{���z��c���]/�jN�>�Q�)*@���	�54��ϛ�i_��&+D�V�)���GC�y#7>7�{��U�ƕ!8�;���������봇S�{(�#R��۝����������dw���^�|Lrv0�)�~S'���EN�9ϲ�?��m�D�NV��<�ˬ33nM��=��=�T�c�%��@U�
���]�s1�Ţ�C�*B����M��� ���g��{j:���!�F�F1qi0,389�HNR���h��j~̙��KF���Gm-����+���fX�f��q�h�^p������z|����=_�Xw3��a�Y�r������ש-5,ϩB�?<�F����B�߶P4*�6dsm��(Sʰ���j�M����&��W�����ONO�3�!��0�|d����G���63�Lܒ�'�VPR��ad/���R���b>
���}���E��|�/vvv�L��A".�HT���@��Q�d���=��-AFA��$�^C��lۢT��W�j�>�ݯ��<�+��|w��=]�n��w����Uw���{� �WAYc��������^��ا���L�C7*[D_`~�\��4
��]��/���]s@l�d͐�J��9Β$�����h�e�r��ae�6����)^���%��Y��� ���	�%UN���e�T7�Tj5	+��np���)J ��t������ϝ���2Q��e��+'�}���?��*�};�k��>@�������L,��xB��?NNN���P�\�Į�������[2��Έ�ŧ��J��M�����i�(�0�Z�؝�'#�pGx���MeBR��im�F���_�.��=�w�YΔ�%.�mT�
;�j��3��Eb���Ok�o�&�gx��H]⏊���_�i�(%��M��Aڜ�]�++���/�J��U���l����o����Y\]�������%�R518(')}FA���&H���Cu�����]���No��U�j��f��+���Ci*ՉfH��������Yy�3�z�Z`>Q���.aW�!2P�����UD���&Bd8�	����G=����O&3�N�9u�Ba�os�񡔈E�؄�جtzi�rCڻ9���8H�&��2����?݇r'�C�=�Lꥫ�F�P5g���mh~�Q��F�_��*��.22�a���t�{��-qf\�	�@q
C#�z
%�U08�E���hbb���
���l���Ҿ��K[f���g��!��ʛ�	N��sHh(�����Dc�ؖ�疖 ���p���200�q��K*�;wºh{ʺ9x�ًf��R���2$:����t�N�s��nꂍ�d�+�=��Z^^�Ж�7�L�v�����ڡm�_K��'L�@�WH][���7@
i� �����Q75�~�"􏼼��w�Q�RҊ���?Ȓ������IG��,����9�m�	'�J�v~aa��p �r>x (�Y��װ���?Ҿ�l���ʌ���Χ��bc_����YZV8jr6�n;���?�]����b���b>=|_Ⱥ�$!�q$�䘫a��ZRFbH�z���v
$d�GXb���F����҆Dm|AT���=��L[	rW�����e/�e�PWǫ�$0�V/��K;�v	]�܍ �������YՔ 8��Yݢ�G8���Ofm���?E�R0��Yg+��Y��X[3 �!��B�>��0N�)ۮ���t�"�n��ϜΟ?��K��[�>e!�բ��� K�=��(��R2²���GM���-9~H�}ɹ]tX������+����-d-e?���=���a�D���}xd��y�䙁W��#44R*�(�u-2i
� W|=�d��k}N�p�@�q���P�"Pec��+�k(���� �MG<��Ы&Q��j d�Jlm�]����O���$�z��5�J�����}|�s�r��#�+��,m�Pʈ	���}#k*I��v:��B%��j�Z��VO]cp����R�;�x�S�m���_���{*66L`Xݿ9�,��iiʅ���Z�\��éIY�G�T�1���#�{Yse?�!����p�p�����kt4U�U@�ঊԢB3;�^��Ը��(a?Uv�/Y�0m�`U�1����KP����?����X�m�%~NʎCSK+�5ȍζ`����޻
�
�b� ���+�E��k��]<��h1�V�����Ё�A�R������`��/%�2�.�#fhHi�x7lV���GQ�%���!'�?���r��j�z+嘵p��2|k��Y�I��bX>�x]/�����  "���5���`�	T3��2�?j��`%�l�
�+�7]~P�_��j�-�������ޮg�N�H�S�6�W��!���m�~{���w)8�[Yoj�>�ӵ�BN�a�CP�������BϘи;`Q���9X/>�Š:�������Z��D�ժ9+ދ	W�X�51666��R���.Ʋ�Hg�g��ӽ=fM��#a�P��5�(�v7��j����T����aJ�ӽ}�z��w���bӣ�Hpz��xy�9�}J��!��0����@��Ϥ>���[�> 	�g#ư�r���� q
kE >�k�RUtz}�ǹ��hB���_~�rs���l��095EE%��2�>��
����Ҳ��XOꃙO��/j�������˩��߿�i��渃W�NrsЧ����\Z=缳R$}��f=����5��MgJTo�b�(����7�	��������9��5�����5vb�j�y��D�����Я�X��!�v;*���o�YY`�C��:�D�$��$&J7x޾۲���i�3ve	��較�a/P��2)��ř�aZ�6�3�����xɧ�p��՘Eu�������_�8;;���^r?����R.U���J�������Ҫ;�6��. �syg��|,�5Ǔ���]\���0���"0DL�W���O�����ՍQ���ݝ��ό�H�e:MAp�����I��=ڣ���ц{s~yO`؊�x�������h���{�(���k�@�$�����fp����f@Tƻ҃Ȇ4����cD��j��{]�D���I��f��k� v�p� �]�!��A����h��5_v捇T�}����D/�7\������3�u+�xl$�M���Ҏ?�}�VYE-�F>�%d��9A�t����#?	(����Ȉ(��-)Q�eX�#������At�N�&���%��� y���aœWY��3OH�8��(����qg䨟_��s5h� �T_�m��|�5t�1O�*��F�\-Z����������))���Kl�ث��EL��S%�j�-�g��2=�yy�3�}>(��р+T� ��-w��4����9��/6+V�����r�U����I?���˘�ט���\�ܿK����_��'1�y�u� �2 0�	I��/�W]�~'2�(�BVn�l7�����F$�;$*�Zޚ�)ޫW�|IF�a1�e!m�ٖ������!�,9�Pc�]`B�~6�k��4�ZҮ�����1�(���*���2� �Ir�یw�ƾ���I��CZ����q|�0�b!th��PX�p�
�ňA<Gp���?�?zeywO�k`k;�t�L�f	.Aj���ӧO8@Y%�Ѧ,(*/���R��d���"�NcȰ���`�����Zc2��rS8�n�����rc�E�j�aUx�����n�D,�`�@P��R���
%6�+��Em�w��|�����,�(;ؽ�"=��Y�&?�1����Sm�x
�;8�/z�����D�P��-���L��ժ����HQ^AU^�L��f�x�2������Ƈ��9|L�h� �Bz�&���]�b����ra�1��μF������q����$��  ���N�i�ۥ�軄vvyo���%m!�pxHc�ڌ�n�
��5J[�ǧ��wB�V+�}� I�1-��XFqj�5����/�mm���e��A��u���'q��yCz�����!�`��ZZ ���O&[�=ȗ*X���0�!ȧ��IfZ�{I�7yK��h�3��(`��x��<��[9��p��J��,������H?�())�x��T�;&E�'Ue�ɫ+N��iѮC ,fy��� <��R��#��{�}X����Z�gx�G�u�e�o϶��I1���t跋� VK�G��`�j�'o��[KOز��H�c6Č�� T� .!�Yr&r �-߼�X�|0o4g��D�������QOj6��e�z���<��&C<��Ci��`���!]��8�G�������*z���Vz 2 a��o�����)��:��I`�1�rTUŖ{CSl������1Z,%���|��i�/�pn���� {��2�ˮ�N��}6�K%@R7i�_�����U�]C�"%Y<q�~h�uu�����6��Fn�5�&��tpXmmϽ�b�+~�C���8����� Z�3n����K�.T�l
�l�&p�*ؿi�뀺����t\�8gT��
;4�j�I~�wLP-$2�����MޕZ����:,�i��tw#!�R���  K� �]� ��-� ��"! ]���}����������g眙��{��.l5pC���\�T�B��]�I����6�m�t�LK�1u����-so����>�X�����=iH@ ��5Œ����1:&́~� C�T���0i).3P�2lăp��iA�sEx ҁ^;v|��Ȱ���p'G,�~�[�NS��������yDooC�������F^Ak�tG��$�$AhD����\����m��)<0�A�iFΗ��7�x�>�.�]���W�%%'G��HL�`��8������D�*�8��J;�P�t����&A�s-���(�1�Vt,�R�Ғ'Xi� ��_�A��˃���e$�9��<r1IH�z��Y��ܨ.M�Sz_z|X�mU6���
�&������z��Y�puI�3S"�a���O!;.`���W�h�����!033���:V��K�������=)*, �����J�}�taƂ;�WV"6ʲ�f&���V�#�?u��^�#���P7+��=�C�p9u�3g�ߒWZp���C�ݞ�����'�=�V �ɑ��S҇@Q11�����@n�$	Xx;��6���1vs}��@Qi���`���䠟Q�-���P���
�	���j��"�����r�Og�|!,:��+1IR-r�A�(  ��4R.�W+�d.g@�)o.W���r6Q:6 \��HHH��٠���͝�v��&\DX�@;�����ȡ�փQ,���u4�|888��-��q!?�c���uNA�����*X{)��@�v��n�X%8p��i�k�*DC!�M��ʠ&U#_q���8:��Y��Zw5�����"�eV��<�xO��=~w���c�(���ӯ|2�uAX%;114rU�{��۴a�ݒY����>���gl\�;_��Jvy}d� \��W�Ø������`��
�7x�����,_{��@����t�bL0�l������19���:�{��uf	tѨ<���|�'�9�Ӿg��[b�$)^!` ��HeeQ�In�㑒�s���O㻇|$�mmߛ���k#`�o�"������/��`��f�t�
���O���:����	��ġ<BBa��ּ��#�#�<�e�8xQ��ֳi����q�ܼ)�3����� �)&߮���hK4'�ۤ$m�}%징-�R�p���Ȁy���·T�[s���dQ�m�O	�G�	��x��D݋w/�Bl�<Ľԋ\�@	�*f�����ꚭ�`Uq�#��V�L��S�w��Y�`��P�u�G�>iS��9��M��zc�#[ �je�W�Z�6���*����C��{;fοo�lǦ�J�1n�����q�����"���s!v�����3+���	����ef޾�i�.@)0��L6��.e.�k��
s�2B'F+_6��u^Y����Kp�I�@t*-���Z�玥�ѽ����r��� ,��e�<5� �M�e�x~q�c��C����Ӂ,���]w�/K�u| �"!���u���w�x12���`�R��U���5C \��j�h�Bs�t	T;��Z1�v�7E�Yq�L=泷o�>�gI�ܜ��zG�ɘ]��B���m���Բr��O��!( >�P:=�ӟ8J	�_���`!��,uY,�x`�0��D��X��i�B���+������r�2�3kۏ�P�
ݬ
Dd�5j����"]9[�22~�bS�Ҫ*�i�1��y&�g�Qd�6�%�Q1Df$�������Tb�E�Z6�z ��4leG��B"G~矎P2��,�GNf���3��j��l�)H�L�EE�Nw���O� ���z찾^ɳ5�$:zzDҨ��7���щ+��I��l��8M��z��žW�������ES"�_��u�ML�n ����s wk�7�5��f���
"__�%;�x������1h~U73>iM���>ln,���8��W�~M�Q�n;�	á�N �t�n巾˅�Ͻ�"��݁f�v��ϯ�����&��8�kyF�13UBrrhB{i�M!��N��au� �bʢy�ZR�S���������H�����ӕ������8$-��Im�İ������F��$��w>7*�+{��靊�7S��<�?4R>).����VB4[�P����m#U����ߛ���hh hj�e��#��dx�P�jD� ��,&O�р:����;E�-}�����s\�J�G�*>�5hu;!;��aD��C-{�Z�##QԾ�%f�	���/JH��%B��z�qq���4(���B$�϶�E�X�g$�lˎ�t�@gNdĠ��$m��jn�)�:W�e`͂�0[�z����q��r*js��u�^^D��o��m}SÏ�q�Pb�z��zK;;rT>�1������?�|7�:'8���D��87�؟������-��;W�.�ʯyo����A�s#����V{�GԋE3:�XR�'�lb7Ic���ٱDu�&����E�3��UT �$)9�@$������T�	g��L�`܄A�[Xn�+���p��.�mG)++3�<>i]� �<6�7L�h��B��������7�ӑGӋ�����u>O
4O�ՠ���$V�$�R�~�K������(�c�.����*�O����ܵ �C�p׭�� �/g��|4�s����e�i6W�V�)G�m{R���V304Ӵ~����~����>��v��SAO�?,�HU -U��E/Iu��i�x$�JA������j>>���g
x���_|��5
F�FA�l�-�7C���ݞ�T������U�6�P�
�lǠ&�8߇���R>|�?��6YS�%�m"�j�hGBڐq�E����V�OGG���>���͐�j����rMM|3s�W���f�4����Gn+��sm�e2��m|���ͽ�I��͛��B��i.c����N��~ ��@�JQb��ҡ��U���3�+CC@9sw:gt�Y9�5>1�>M��u��)��������I��`�
�L��������9
D܇���j�O��ж�/��z�!�3�w�H3� ���\��.���j(��M?FbzT^�����o������� ��4�,tqqћ����j�Z(hV�u��p/^m��>Ԙ������WP��[Ӑ%>8:��ʘ��;Q�>wզ[��+H+?��P�����ZI� 2"Ӏ_�Zhz��[�%�۬��ϭO�=��n��!�[ C[��q:�:飖@��fHK��V]}�]T���iE���Uk&ĥ��-#��.u|d`��/_l�3�I�`v{Z��쏀�D�5���:�ov�ohh@ ]�����p[dT�މ�����.��>��5�;�d)�|�ޅ�����{���js�f"�=:#�b(ݎ�ףa�t�����iiRVr!��[b(�H&ʅ���9��8����*.�R�[���q������Y[�ks���t{s#Үx&�Q���Y�X?rpP>�� 7'��
�5 �W<�Ү���4�$������^]]9��h�]��U�z�(y�>�yO����Zv��ڼ)�{��@�E�b:��t�u�?�}�P�L��/�N?����և�ys���1U[�_B6�[�������l���a`l�?���2p,|mK��D���+��:�ŗG��������bD��.�^�����J�QQ>��F�ӕ�4�h��<>���bMEY���ʿ��t��^ThONO�X��&ྺ��[����d��o���U%�1�7��~KZdɋ/�����%�B��߳�|��k�9e�ФSk�V\��@%�o:D��a��(�伟
KG�c���C�,g>6�\�#7����B]n`��V�nOhϿҼf"U��	�s�&S�b^G��� �|~%e��J�"�󴩰��w����9C�d<��3I��K'�5q�/�9�<��� ~���}1w��I:��i�����VXD�&y�]�c �Q�c~�Kp���&vv�F����Lб$Ʀ/����б�d��a�{����䳾� 8��R�F��E�n� fi��͗��e���a�o��++���R����Uؓ�zo$LT�5�؝Wu�Q�y�U��=��!$($��Ё]%K<
���^A��0���X��377gJ����9
gb�;�B%�JP0��Jց|YHCǃWPPл������a�<��5�Z/�RRBW|v6l��h����L�y i5d-�G=M��9#d�2@;/��L ��ʺ��_��skJ���3�eI)s8I��kg��4z���6��ĸ�kK��A;_eS������O{�f�-\Z�e�j�°^ZkR��Kٯ$jdI1b�ć��}.�v��{���k���%xW��~U�M�ѱ�����Vc��U���<��'�:F�J���K��F@
8����S��e$ ݪ<"|��s�H2�~	n�w��1%��c��:3��=����V�ڗ��?��Z�a�'���e�?S�Vx�X��ojJ���:v-lt*"�K�Ƕ�!�Q��Ї�St�_Y�~�i5e�pZ�-^n�]�O�KKK�Y�9��7�6~���S���Pg���p>V���I�i=��4e���r�����` �uv�d��<���D�f�.kqe�SOO��*��g [z�Q!���hM�d��W�'l��'������h�t�-D�LL��nE�/�vb�.P��D߻'W�����'�UO z�ܜ<��HA��v�-�>�e&��u�-,�LWԝA�%o���`�w~�--N���Z��V&v�R��|�	ʿ'��9u\n{�v^H呺dr������eZ��s^z,�
={�u���rz���1����;>l�d p��?�8HJJ~kv������W�	j� ���
ǢS����ݷ���}H��95hܺY3.��Qґ1mB�B`W���=6�x��eA����.#)��ݨ=З���OCCä�D'F��7�C�@�S4p�����/���_|ϐ%i�FR1#���M�v�E�\d���wQ�8���wF�3��%=l����k:>����oj"����@��@��%�{9>/���c����X�|U}��-`����WW�o(�����㔝/'_���bL���:ֈGm���G+��9��M܂�0pu��)����r����|�DF�"�믦��>��3O�2pت��|����"vKh�f���]���[������m(����F[F�u*���6>K��9'15`̺��(��d��;��V, d��w4r��	D��y/̃�
4}
tYE1�Y��J.5�]�����5�|����/0�噦���6oЇrP'�Co=�ku�N�K�&�k�ZG+����)�a�D���/���G��r���Ͽ]������zP���Xh�힞&��h������ԣ���_�)l���6��aK3�8��kH�Ǻ��?U�o"�����,hz7��>�	+!��z�憥�|���>22�S~ENdlp0�����?�T�?��և��F�!F���������v偓����k|��l�����.;�f'wB�3HBB�^AO�W>��c3d�X)�������@Q��N�~*����+Y^���`ұ�3d\q֏.��z�ml�<�ng�76�q�g�����6�ڀ��}�(,�?C�;s"��f	y˒�#,�w���E�9P�ց��P����������9Fb�sfV�)?��e����}%�*�Zj���	Nnnn��i��'T�dI� [P,�}����h:��]�<��:���Eڛw?��t6�<E)-\��ۧa���q��$�T��2�|2���/��mhpDF��ü����oّ건)��se#j�}	�G�+��=*mM���' [�W��踧Ǹ���M�� ,0�z�d���)Qqy	4�)�_�ŋŻF����*d�����A�솿��7��\^�X��_��9V���z�H�v�"�� �Og��2��)(d��1�pp�M�((0�t�+�!QP`���RcF?sXTV��JN��-��?�H5������ �l�A$?�����^GT-Q��+���"�ˇɄ�T]�Ѵ=��Kn�� C�m;���Ѩ�? � f>@��iD�[f]�zj� �#���u�s��h	wK�7�9�bS	b	ٞ�$s�%}�B]ZF���+�#;�u�����)N����C�&E`
��܏����RC�?�7�b����7��U�J�L!�/,���઩)������y�D[��z�����y�.��>0���u��AC�K�Q��X�_3���P3
���.�(�E��Z�#�|4G��B�����d��@FD|C�|�es4]��|�>������b��YғZS�Va�����`���X�G�i55\�ëG�W�@诨`öz	�k�e@��q�=���cWXa2!;�v����E���1R��+Im��7���k���� D�2	��~}�'Iyt?�̔4�w�>�HA��f����t��W ��y	���I�8���a͠�m�E�ܵ�i\�f{~�����h��#i���G�F����?�9d�H!���vRgy2q�3_�廽���usmu>��}�RZVj�/;�}����9�ڳ3�4��}g°��h�F����hC�hYʟP12*n��
���N6,;i�LO4j��%z�R$=+^/�����Z���l�ůƥ�Xx�ɍ�yCz�ZQ[�6�o;���LE���;삣`%��z��G!=�p�t||��>�.�D����vp�n`��B��	��y"c��{�ϖ2=O.S'5�?�ۜ9s���w�\P���Ll�;�,N�����\�?v�9C����̔�KM2(ٽc�Ar��ڰ��_�ϯ4,>��� ���2�wr�|�q�F�f-m�-ETttn~3�rT�"  �^T4lwn~�B�5�Ji$IG�^�щ�v��_z������ȎI܉ַ�WeU�hr��}CU�mP}T�Ii�����zS�00ԫV�y"��i��u����1����=�q;=���ցtba��'E)�wN�.�-���<{n����a7h���3���b1��q5�t�#.x_�Ue)��5�2T��(�x��sr�@�#��ĳ��O��=ۭLL@0�?+��d�#�z}]cf�Q_ϻ+R�h�@�4��Y�h�p�]e59�3��_3�}vI�PHI�Ct�޹���dc��1�t�)�)��T6�;W;�U+�?�Ɂ�A�>��3�HHgc�T_/O���t�P���Tat'G
��J�먩�c���h"���(�ᨱ�N�{�����=3k��A(��_�#f1�4���=o�z��a=2��=��rf��d��J0u_VN��X�mqq1bK�{�^���U���/;��ߜ����9�=���h�R(->���f�~ �LL-�*�����!]L�c����=s�� ��B���5Y�m��ݹαxǴ�Ð��̏�e�x_��P/x��zy�l2�F) �u��V�?k��.�����)���;�o+��iOC���h?�q\jX�~���1����qp�ц��a�������O�1���}p�����`���Y�'V�������/6���eQ����z�e����1��j�>�6l�0���=���!X�̵�>�2S�3wq�eT��MG���vX)T��z~�W �*1�S��To2��ml��]���cx�.;������hn�(�W]/p�Cѷ�+r�J��:��5߸[]�i}�욒0O)�:t��v����(��ag�f/��5W�k̝�3s��'�	X��|�<)���B��b.�%���r�R㜰0��0���6^T���Y����f�3��5{�O����l!=���g"�ʴâ�l����?M��芟춍�mGek�+!�@�s�PL�v��,����a��^a�Ye_oo `�����ZJJ�5b^W��U�!�u�:�=gӕaѴ�S6�ZZ��s��ceG���H�pv���/3*����q��N�M[OЭ��jxH�B%}4X�=.nM��w�Էp�(m����T%k�� �m�ש�(��A<Y��;�RJZ� �hjjRss�� &e�ա��酧��{����g/�9�q�$&'���}�Ȭ�j�n��>?��$��?1��/�
/kh�WQ���1
G�Ni��W������V�`2:[b�-9&�"Vb�AWC��Zܰ�0��Y/��y8-�lHHH2r8��9mmd6�@�]�=>��z#�|�2�"�$1��}��cICuux3ȵ�33��ñ���5�=R���9�9�<~Շ�	z�uM2tĻp!��6�6A�e}��/12�#éI�ME�`�H�43�`����w�bpu�nƎ���Z�z�M�S-�Wx٨����4*Ex��A����J�W;�;86,�<�[��o4�P�B;��No$��5����YD4��� J)��L-���׋^��rڋ ׊�ܶ�xJ�wF-]�)�,.��䔖Q�cnNV�3?қ��_�M�`.���2h����1���X��9���p4+�iT��R�f>f�l�x��Ș����U's��9?����]ZU����6�fu�Y�*X���� ���b��=�=6��/,DH��y	��/>q`����٭��gߘ�gpc���� �������Uб"r��%�1���0 ���#Q���������"�dG@C# q���_��
��&պd.�o@=$�����w�����S(`���3u�t7��o��9�b��.j��x��EG�����qqsÞ����)��$�W����r�
�RG'�)L
�?��#�����kpƮ]���\||�]o�Ǳ���� C%nm���B5��_���}�gR��?BXw[`�-AL�-�<�

�/ƇZ����4�����0 ԹI�f�yؒK]KHL�'��Cz�Yt�p���Sn>��%^�Y#g�0k��� ��QYK�A3�͇�.����Ѵh<X��lh� �����G݈}w#�M�j�&'y�Z4�c�2��(����l
5 Ҙ�NF��ϟ��)��fa�%!!����6?�k�2�3��gg������^�0U�z/�C�g'�=ݗr��TPa���ϑ� �������ϒ^�w��os�ܥ��I����/(�Mi8"gHx(�7�<
Y�y2!=�B���VY5�uq?L�KKc���p$jYG��K>��L�<���Q������ ����sU���1��6��>��_�{zz�l�j�����ojZi���ܵO0��n�F���v�^w�r�k˕V�^01���:W��[��N�[*⨧%cf[��D_�ʯ\L>	��OTdj��~�p��
��&$�F������r��@)�|}��z��By�_���d���]� �mK.!>�$��M--ӹF{4
9����λ�Wv��r�x��ͬ��K^e���udwP]�og���: |W�@"�j�x���%�Zs���_d p�=wE@\<������UX�� 9�k�XX�///g;HۜŅO��|%&7o���pȹA�}��a�#��B�J�2��P�FX�����xZ���*)�| ����Π������q����)[]�'9�}A��s?��GYHyxL�������@~8ec�n	�cn����EI*)En
�,7�jfb��5��R`0�g
��6w�-����5��,�]���q������P��Y�8�����V���":&&yW���ui>R���G=EG�� = �}��e�ʁ�����%��o�D��ߵ>*���ŕ٠�M�i�K�	����7�h֔��c�`'sL�Koف؎�bV���?F,�U�8,��	2ZAg��
�˂��9<�b��E���KB�C���\~�}�ד�A�����v�@�.�$�-�(�6�A�\�����|���]h(
�+�n�g�S�\`�s��z9�g~g(b�N���ָ��
@ƒ�m���I�q��8]e�tE�==��?n%feQ-���4iS�f4��n�{��+*B�E���>�Ӵt3s���яFL�\����U�T
���h~y?�Aܟ�.d��\�ejЧ��;)E=���@���o~DJ6�����~��'ަ(?�As�+�r��k0�������Cσ%�w�����4��p5�<���Z��=�����ꮛ�	II�kb���2>��3*|�)���I��� ��p��[�����?\_|���6��_%x)Ȫ�TJ���?PK   x��X?�-�,�  )�  /   images/6217b039-096c-42ca-9a04-ba011aa6a0cd.png�PS[�6*ҫT�%�AE������&U��Հ �"HWi"H�U���R#���D=�|�?w��ܹ3w'���Zo}��]km�+J��;w�X*�|�&�ܹ�x8�7�����&��9)�?��� �΁��H@T��+��P>,� .�oW+���Q���v'��+���˜w�P�	_��ý���g^y�m�,���
��X�ŕ�W�0���q�#׷�f�]qM�.��qPR�Tٗu����K�[����frI�<�����,��F�f���W����S�I8B������&�����9�F��\7�k7�uW{�6�v�B�i������� ��ŗQz�s��L�P׍�j�/(#7����h��`����������'�S<�����~yndce\<��_�٣����A��3�tA
�5E6�DvzɎ��pz��3�%��!>����I���
i�y�]�����x�p��+u��LU`;~�����\]�*V�&������g��D�k��4"Ϋ[�G�O�5��_R����U�ڿ���Qr5}u�[�蕬gr�4Ӡ�f�zT2)��_��:%�E��`S������4��	��if��]�I~�W.�x���IK�ָ��
�L�I��j0F a�"�Xj?�������2��w�S�xv�^焮U�p�O�P�<yvK�i��r�|t����O^���q�g�p?�P������|=^�H��p8�IK��m�WPp$r����԰�L��80,�透gB������ӟ7�o#G(�8��B�V�?q�����9w�����y_�/l��%S}�����E��52�����::4�t�;B߉�.�`Tt`�*���ѝI`�p����-�:��"Lw�q�<��v�] �����/���Js=	�OdZo��ʴʜ>�������`�K���w]>��d�/�V�����" �_�E��:v��q{Na�	�PVA*N�+`�x�iS�8鈃4W�?��yy�V� �j�Sc�f kcfGV߯���joaޠ]�/p�s�Wk��<����L��j��!U�ҵr�{&��+�x�
@q~�io����Ν]�7%!�����D
��L����L *F�����bEڈ��NT�p	����f9%u!>"��gӢ1��E����b����}i�2.ޱ�0�тİ~���s{oP'%�{�VZn��)PG��c�g�A޿ 3s/b@y&��.iT5b��} x\:��4v82��4�ls���bLRp;ݱ�a�N�Cja�6��!��,V�b��s��-�(e�m�J�n�v�6�'o��
"��͒�4��q����,�Op�e&��<�ϟ�4r��� �<�>s�����hun{�=������p���]��J�Qw�0����8�$K߫�u1�mmˤ+���GQ���KЀTGŭ4��#t���6����*��B}�����	��P�G�
�����*���ټ��-��:�+ZNhn�������|wrXs侙@ü�t���>�?d��;�`v]a�G-��y5���S�j���cB�7�3� 3p�(����ɩ�y5��@��x7�-�\�v��hT���.(q���pls�h/�8��7��Paë���� h]��y�M��>���&��>�T�i���Q#��[�6ҙC.D ����/!0-@�tO�"��WO��4�\���n��2��1��:���d��.
^	���b�%l曤nP{o$c�`�o�@�����<����-w�E���E�	 z��}T�ܼj���+�}*�S��T.|��x*#�hLgP�)���i�l�_�g�������1�feL��W�O��ƧD;��9ǡ%����(A�@uLT?ϳ(�b�;�3����F�q�(T��=�rj�����]�y׶#Y������j�
�aK���-��'pI��Tx�wU�@-� ���0�a7�Ă
�")`��7�P���
��UM��#q��.�V?�B�}��q��r)g��Ų�tK�?�e�NȦ��l��PQ�.]c�ٰk�ؖ�°�����p��1�q��;U���:��nlK#���@�ݍc �l��$t�&Xc)�(t �$�S%>�q]�8�r8a�mކɨ��7w��C�PL��{�[�Ժɸ�Lո�Z��!�$�yXE�@�D��^�j�Z
�f>3Н�e]I��推�)i9��|]T�Sp����Pe��yq�mMja��������ZF�A�ˆ��#����[zUI����N�/���7a�!��C����=!)����Qe��4_�1��&!�o��>���F|T�����A�_�ny�,ͅ�����4h!=�W�f&��@���J?�7EP�i���wB�87g��N��\����.#0�m� �dH�J��f>�%�u٨+�T]oT�rR�5�e��a��&����g�3��v����=�|8en��s�ŸE��6�_A����cX��}�;{BFpʶܪx�>��[B9,}|K��g�'3>��33ѡ���,�q�m>AAT��f/�^�Rڋjӂ��ޢ�������$2nL�����vP��K�R����F�� �M�@#�ƱqI����i��E��֚њQ���_�!@��\�Q��c-|A��}ef+������s��l�(���kǸH���!���(J��R��E]8�X1����>��0�6GLx� J����7�N�?�|�T�f����0?Thp�='�]�c0�ҒT�����sooPҜK�����bX�^43-[IK�$k�ߍ�l`p���o���g-
��Wy��7�n��w��6M�����bZ�2�t���8�wc��Pk?h�/-`����s�_j=�������r�P�H4����V��}���h��潙o�ב��$��}9��}�_[��+l�g&�{n�)Qn]�!6��e�*�sZV������S�E�Y�j��ZZ��[>�6��1q~���N��n����*�*����p�pZY�^b�WP6��a���=0� �Fa�,γR8->IIK/i,���_b�)n�4���� h�����\�|�-I��n���+��=�!�i�ɘ�UͶ\�'���M�����F�T�u�L��Fn���Z0;�L�,���/z�jZ2϶Pl��[IFOO��jo����Y6hq�y�a@����Ĝ���o��|���Q�ɗh�L�J�_�'���?&;�wR����Z���ӑ�.ó����	�C[B���[v��R�`�jRq�Nѩ�) �����k�����0��]������1�+�NKMs�L�Jb;Iy�ůi{�'	�l�X�*�f^�I� �o���_����pޑD�U�|�7���׽\��t�K�4x�9�U���G+�����Az�c��๤C*�X��(y���M�v�HcSՎ�G9_�Łt�2�u9?Rx�|�Q�������"`�$�p�31N�Z���rȏ6wk�(���e���A)���sρ*�ն7�h~}�wW��iZ2s��&�?G�;��3��KE���9,�Q��|w�9�w+���a@��8��r�CQ�p�SC�C���h.�X�Ě�L� ��X4����{���}<�;�C���9'J�2 4(�����dA��?�ȃ��	�,=����7J~����ǘ�����=��>!�S�-���<�1�J����`�0Yr���e� �p���a��';9����U�N$[�9e�ZG�r�/]���h��L�X���E�t�O;��]\;:m�v52�9C#J!����`��a\iB��u��`���I�'F��5d�l�t��&�a�Q�b�}���O���-�
�l���}�ד�	ȍ$?��S$1:X��ZT;�J�Q�Y$�D���a�;���VҘ���������< {l��z�j7���t�.6�\����:>���|Y�G
0�|f S	�
�� ��?�k�������C��D �������t���߂8Ir�丳[Uq���PDxY�����P���a�^��l���fPK�-��ٕ{yy��a��,�������A�� nf�4�����f�Q�P��7-�^P��r�Ե��El�+�'�#F>7"���9��=B�&�Kfv6��ȴ����ω9���o�܄IЕ�>NrO8N����J���;�>im��l���7}�,XK�ҫW9�~��2��Fl�f�8�*]�Y��C3��E=^C���#1�ȫl��X4imi�R���OF0�p��co��Lm���Y��`�O�|�d��:�{�"7����y=6̱���bߵ��X�OO��l�;nҶ)��N����ּ�)njm�fo�.�lv�Θ�m�X0݄�bsRP�	6��e@�q<3�n��<�	��N_�[��J?x��x���l�:6����k�h�-�Ī�T���`��}E_����O����3	��^<i��Q�t+Z��6��:�>
���*��K�7C]�zS�����%^��M��@���Fz˼}�x��'?���A&�ȣ�ߙ�x�^L !5���b7��B�45���s�F���X����'�G X��FNk w?VtԿ���|�OIS�COs�].�*�csHm�h�U�6�W�O�?��l��Nڭލ�̷.	����<-�m�߳��m��@r�|Cϟ��&@�p�	�`�^��t�8��ɏ�����eɭ�qS����Bw�Vҙ)b�F�;�R.��Vg���jk����il]��dT��%$����'5��>���<��s�R�Ey�L�-	/��A�������66K��k��`c''&W�L>"3��B߽�h>�5���m����ѭ�U���B}�.Bj0iق��W7��w���R��$��l	mX�"P��7��d<�i�BJi�R����K"o��������ī�Fuw�3�oDn���o*��DfZ!���R�.���<�����7!���vO���&W�R4-�MuiTha��FY�^lݹ���9�������dTҕY��G�[��١�����om��f*���:��>��@`��8�gu����bT5�b�i;2���9:{څRK�����y��?9<j�ޫ6'm�s�2Bj���K<�����_����~#�=�H3rzf�~f�Ѻw����	�N�5��m�E0�<W�N�S:�^}�Z�Y��"^X���>�"h��&lJ��)F�=��g�t�T��X���[˃�ѵB�z��h��x���=Br��j9�����#�c}W��,]bEz
�c�9G'���h׾�j�U��*cl��h�s���OMd]bu�*��Ɓ��Ǎ�;����b[��W\����K���7C�.��]���	D��t�5BM,��������6����1��[�c6��=����hA�M�����D�U�#��D�Uɦ�u�T���2$�	���R�ZQ�E1\.m�0C\�+�Җ���0��'��op�gNVW��d��@N�
i�w"�.��F�� 	�������g�{Еż�-#9)����LmtQ�IG��]Ya��")4G����
?�{���#����#lH5�5�y�Nî��-�
�u-ݠ���9^��|d�~>�� �r8y����s��/Ά���(��V�����m0p"&V@Y�<�x���}<�6�w�uB4�.f�4v�x��k��W8Bŀ��z�`g},E�V�������O������?������OUh왵�b�|�7��T��1�82�$��?��@P�����I�{��wfܠ?u/���-\h��}KLB�w'�]��ڠ���;��.�}5��K��{��R��Mwf4,��."~����W`Ц� huE������GI]%��@-��Ċ��Oi��mH���,;���^t�8�s�h��첿Ŗ�"~h ����f�&���|��H,�7 h@��l���2W���c��R���sl~�����
�8ek�ub���\Ɲ�����M��X�{Ɖv(�|)�<�x_F_O�9��z�����v�� ���\A���&����ɢ��(�{ù�g������ �q9'����?j�Ō	�u�c�?;n����g4�# �����j��;7R)B�H�&!֗���7�� cA�� OPC\+�G�6��mZ\�2�8.�����wt��[�Z�w���ìͻ-R�_Sk��|<L=lp�j����`��ߣ&Q�$��rynY�m�Hjet��+�����H�#��G��"[ǔu�<�p�~�l�����"�;D{�!��)O�l��喷�-�V�z���ŋ���v8�v������`��0�ʠTe�g���v�+�ս�OD윌��
��*P쀴�$jZh�/��v�lD�m��_g8ev�f�'��x^�ܰ�:S�b/t�Z�I&��\�r��85���^@��;W�{΀��	O�6�|�oþ�Fx6�P�kVcW�������KR#>u��{�����
e*�Fo;���v2���~7�	�|��S#��9=t����� n�7�'���?��;.g�yL��מ����d���PR-�:���ލ:BϤRV�q\�ܩ��C%�R�	�Nŭ�,��-��pT�O<DK���- d������*�\@U�9��78������������o��}D��D�V:�y���H�mA�'G�Qw�E���}b��b���q]�b�����F����t�������=�N�{�o��+�m7U���S�U�B���������������v�?�;����c (�a�����������9.��iܓ�UUcΩ�k�����0��d����
�.L�
Ctyp��<�:�p�v�w����g����qk$��/Q�țk\ݺ<ƴ-`g�>�W�@��~�)����f&���m���c5q�Y7Q��Z�|H�Q�|M�F��<���Mu���G�r`�o�}�׋��tX����T��E����h.�!6��6���3[�qC�vS�p�G�t�g����%D)é��0�Y����Y�������@<�?���B���Ld�+����,H.y�7�B����e�f�}�����#��q�� �fF��| �'�iՍ~SN�l@�n,��H9do��K�ɹ�,>L��ȟ��-�-�idD6X� X2^D��H�m9T�:����i�]�w�69�$�� wm<�" 0����CtRb����:�{w˃DLZ1��I�CM�~K��&������Y�c�[T6�]��=/��b�^�\@���ϓPx��w]`-�����t!�?&������D���[��9{RK(��-��Y���d:�jf���_8zu�9, ��,|��?���dB2.���w?�~=��MĦ��}=/=�����%OK��݈�5��؞�:�?�������Jm���)�vU/Mb�WU+���[��e��D!d?����D���l���s�?֩Qe��3���9�̯�T���"=5./x�q�{V߿8��<mg��٩,u�	w�J�T��YF�Χ��0�[f�]�~7F�� ���Z�A�n#�z�6>�mJ�}����i�O���暕�Yb�?
��Z"բ�����kwUOT�4�[1�y���`8W"Ə�"��\�b0�Z���	�����J��s����1�R&aA�V���cز���E�E�=�Ӈ?�1-+T�/V/��"��"~0.�Us�J��y���cAbT&th{�U���k
^�O~>�\��;�6U&����,s�U�˴rd˭���p̥���0�� ���򵟆�|�Q�e��U$�@���1k8ȣk>��d,.T%2)��|qIq��̝�����������p��9L��*g��
�u\/�wF��?E�4zH
"�����+�������p��&5��f���08�HIO���fW�rXtb�����!�s���R<Sl�)r��A�nA���*�TX\����HW��?��I��^}0����Σ_>�h>Wb��̞c����������G��P��G�"Y���ja��G���1UUg�SN3�u��.n�����wB�!����=�
�������۪#$H��K+�o޼�\���%�(a<^V(#ʶ��Pvx`��^`��]V���R��3�o 0��Ν2緄]�n�l���-g2�*���d�xz�з�O%���Ӳ���݆)O���柿&��|]�0to���p}n+f� Ê�)�.�K�i;��s\�B�;�,l!���A�����Ko\�[��4�X�~���~f�|� \�OXs�B��=��jl��K����� �\ە,_ls兡gT�,�$/�/O��̄��FlP�~E�\��a��@��E��~E�e�ޙ�vO4웣|*�{�������� ���#p�9fUo��B C��x��l��}.h�9���m^?0:��_?�}�m~8C�R�@�RU���@�P�ɗ�Z�lU�'���bJ��m���.Qz���k�� ����g��2}�7�������T��I��`{��
x<|f[nqY*?���
fX�0�UQ�D���g-�hY���VM�-���)�cH1k��_�����/�Ɯ���o�޿}T�Y:w�
b^��'v�gJG�9f�OW��^ 3W�S@��G	��]r�6�J��f́���ъT��}��ۛ�By^^�V`�_�_ab��5�CǴw1�i���z�<���
��?9of����5�( ��Em;wך#8��^���&��Ux^
��m�a��U��9G(�@g��SIF��hn������� z}�z磚�>^	�>Z}"1�k�1SI��q�M�}z��B��v��%���}$�s����?y������F�^}�u娛�e�~:�[m�<���6U+��B7�ri��6���+�Mvg[z�d4�:͔��*�.n�,�?@�{�������1��%��]����l�����͑_�0ð4\.'���=1�0�1��t^e1�-��-������j�V��z�H�(gKO��B�����_�y�����<�������I~�׬�n�O�p?�Y.s������TNw�3�Y��̅Ɂ�����z�7�'����Z�DD�����z��pg��8-v��l�E��뫥pKccK�����,�l�ΊB�9x�/��3��oJ#H��x,x���$���tL��k 6צ����>�;w5$�>P�H�b�Sy��,�Ui\���Ċ���z��xa��-���U���㮥+v���s,�w�{k�ۂ梩��F5it���,B������2��>w�]���R�����u�+W�jQ|\��,nA�\)�P�����r[q�|�m��S.��X"�b%N	n��;��:��G�����V��y��܃sf��Nf��Y�^_y�cŝ�ܯM��:&���n��06�>h����=�c��.���!Z���!�[��y�M�J7��bU���"�R;��������yM���,�2d╵�	�Ȝi?�mϫ�������?+�nX	jWY��3j͹�x.�A�Eځw$��CXp/4~�����5��rp:�M�	N�#�f�z��<�w�ۄ��c���7L��p=��Q�ς�5,'=m �|�˺�+��3-�o����)�[�1wF���$;�
��z�*��FF�+x�x���d ]"�+�/���)�W7$�u��ST�bշ8t�G��f��� �XT�d�t�4�9'�$Bθ�M*4���bx�	mwU�@,E���}�BNe�Lj?��+z�����(_��u�T�ڷXNy���µ�׻lyw��v��pYj����aE�WG��&��ݫ�>��sgFF�K�m�������D:����+,�t~�ݼa��%��I�]{�0�ilk����z�|�`Bt��얫�c�ј��+J�U�z�T��b�2t��p�:!�sϵ��'m���^���$�[��d܌��L;�5d���h�MGo��m���eX��Ӻ�N���&M�e"֦��CV�r��b�6�zjӈpG��zA�z�
��+�)���?��:b��pS5䫃��Q�kf a9�>�k0��X��ȣ1�1P�(��y��ҽ{�����'Ȼ������Q�v�\��{��DKD����'v'�B�-�ݵ�����W�5&xa2Q�ˮ@!���0T��1��6>��46Y���
p�<ˈ��=z�R���,ڕ�{�S��v�r�M�t�~ �Ί�>W�?LS]�&I��\�"Y�]�a꺞�����+R�.��&���<���kd��_�h��OJx|)\�?2Z}�;_�a�"*b�I�!����+�7�����Sz���Хq�e���#�z&��nDw���ݏ��V�axA�0����H�M�ůWY�fY��WJu�S��rqh� nE>�E�<8����j@
Ξ�����6�r��eῖ��!kU �	�E�w��'����C��Cؔ更����W}5ʺ6�.l䵞/���`��\�$�+����a�E�*��>��I�
d�1���-�f���u_}����v���4���B�Zq^k�S&�/p�S4�j��%�t��zo����U�f��+j	T6Q1���D�Ev`q��=yxbM�H�s�F���H�[a+оt|�K.9E^�]l����rՂ�|�M}|ik��o��':�B=��E�W�<�8IN�W���Yhِ�`��&���p��M���rm�e��:@$����Eמ�כ>���c����� `[Oi�^�U���cL�>�;�����FMm=�"K�g���PX�x���_f���\��>Y�]�L�M�f7�`�Y[W䀺�oaT�E��eI�I
ժB�y�C"9�DKYGq���qN��m�D�t®d3n(C%�U
@M1k{*���' ���#�{�j��O��* �fi����:��{�pp���`�ua��ǻcH|:�U��.�u?�����Ȫ�
�^���2W�F�R��?=��q+\�OU���,�=�d	�=qS�7�;����^h�<]���$ɿy�!A4�F\�p�AD��rx���"�7���[��KP%Ú��G�ǫ��Hb@B+W������GeL^]r�[kN��D�&M�X�k~yQ0������	г)#�4yrL�>5�?���c����9����#�{n!ftA*m!u�S�-��X�N�<�A��ʻ���k�ZK۳��?m��J.M=�{++��Y���~����:����.c��2��v>)+-��RG�eV����'ē��y�ה#�٧��b�A����`B#�>*S����O���M����]K�O��b3�BxJ������ڬ��E�"���1f����cO���m��ק�7<��#i����<�߮��������?��>�$���%�(62J�@z9C]*���;�nNMA�~�^�λL�ڇ�a�v?P�E�5TB��/\�:��ד�ں�m�������>`�O��ޠ�{$d`����A�@��u��ev�/i�#v<S���9��o�Yk���_�W����}xWh��4�PD���ȹ?�ir����>;�|P�K����<�x�v���'�B� G�����8��]��H�L��������[%.*#GU��F�)�"s���9O�Q{_Pi?�=#� [@�|��F,i���_Occ5�����־{H#�gC�(a��Ni�Ǳ|tد�(�������<$��b�T^CY�j�U�����C�VĬ�*��/��o�ۓ�GY)�&c)�ub��Y;-+E�t��a�9�����/�����S�b�j"[���U��u�B:?jV���ڞ;6@�6~Z�W�4��a ����j����7��l����rER���[� !\,I�xb@��Zj[+�.�yX"`�Ch�Vd<:D��
��ZR�g�zP��+X��u�D���nf��!�a�7[��?�umo�R9ym�TrPKݑ���'�v�tan4��hw3¥��y㑭�*���Q��(,�J:�� Ʉ������c�ϱ���.��N��3C�>����[���7�[�gp%��YVq��Z�W��MV=�H�*y0�#�'�k�/�����Ī��ozLJ���L4�U!岻뽈��Pd����v��`��=|����*���ꗠ�2�!��m�����d䔵�D/r��A~"��s���^}��j���h�d�� x��Ȼ��y�qhqG|�4��S� ��tY�5���Y[���%���`�,%\x-���]D���`T<rN�i�gr����;�uL߮-d<H��zŲ�_M=��(����I�#�ڮ�6*��st\��x���H��Xsk�T�dJ�R�/�v}.�ͮ����"�kc7��?�E�>6��w�����y��}�ih��_�Q6�斋z_K^����´xʦ��r���B�!��� �աB>ɼ̎��s��]�<�1dA����lO3�H�[/2�b w�&�#�*�����k�g�sCT���OW\s\-�f/`�N9q��ȯ�?��Q���~�ƍ�|_W��y���D�xl#�;��e��|��m�,�l�|k
��)W76�p�����D�j��������B�_\&9�	a���ct2������8蝅��d\9�<N�.	��J �֡��@��\P�6Ч��
^��7C��!�i&����KIH�l��wƸ�i]�,Y�}Cƙ��a�%c4��On�)\��8w�o)� ���j"�*����o��bg5w&�z)�l�W��E�<}��.|L��J�G�M�/�!1�U����}Y��A
�l�T�f��Bw� ������9���?�uz�Ѷ�\s#�R�X��^���G6��I��������)@���(�xP<�\h�����*�~�0�~�`����s���l�k�N�jA���F,	u�2�-d%����6�)�%��eG�;`�Ul��w�z���XS� f�,���nǠ�?o���b�����o��8U�*�S��t_M�ݐ��M�,M P�}p$L=��c�����;s��"�M"�����|1]>~#ao]V(,���eki��+�q�O$�k<qdMK=|"�(.O��tZ�Nr�4�.A�z��B �P����F�f��e�f ŉ?�8ܶ��Nվ�w��{"�r�f/�̚U�=�-4$�@,��k�$p�=2T�{��V���0���奐�����Xa��yS�y}�R��m�s�̢=h��s+:7���@X�7���W��_��9�����q<��{�iֆ��C�AuƷ�����a0��V���\B�;ɻ�	��æ&S/��5����_5`υ�Q��3��.�J�Jt�t��e-���!�����{&}T��{_��dGo�_|w�P�2����O���;�_V�R�[уĨ�BwN��D�V���v��m�;~�xwO����R���)�շ��.f���qſ�e����X�����w2Vӣ�����$;]�:&Ѭx�'�g�v]��-��ݷuaX�p�<�O�ؠ�Ni��+�<>]5̿�٥�4��y���zl�b}o�0���f�oG��.~� 49�܎Y]��6P&��δ����/�!���}I��=w@�Y[[��GG�Fs��B��EW�(�g �C��)�? s�/�h��5pE�a�Zl��G�ω ��Y����
��8�1�0Q78�B�Cj�4����X|�~��5�5��F�&�?9����Ź�a��4�tF�	]6���YX���B�*f�^�!%���E����_A@����nɒ�@@�������
�us�%B$�WT���=��S3L^z��������tM�L��
��j�]�fa�lg��o����nԀ$<��5�]����0�)�����_�U//Z]8�țgnn��4���}L���U^<�'�����U��_'�N	N>�3��}��r/?��ib��8��[��d����І�1�Ƙ�%����͇]�&��!�����@I�]a�&����b�k��=�h����@�M�K-V(�?IS�^��f�	%��/�0�ҡO�2��4�\&i6���>jS��}�Ұ<��L�m����)�\� {ss�����X��LY������$� �!Y�}z<x�R�F�7��EOޯ��+|i,С58h׍�[��L����" 㧇��w���i�n`B����hsOd'R�
+�X���Yh�^��Ymޑ �\������Wu1��N�Q�e#�˶tQv���7z���M=��T��)wWۋ�P�e������+��{�"]�&~�ZE�u��0h�;�K0*�]��1"�B����>$�����#�Nf�~n��O
�p�mZ�e�Py�ΦEi�;���N�ܩw�� C�my`2���tv�tc�td3n�@xM�Õ-�[9JԴC<��)��=娢U&t6}���^<%����@Q/��)�PI�ѝ�l��e$�
�.K�E�Z5����1�@ ��\�yx���RE�x�����ؚ�,�����lB�E��-�m*^`��̟��� Z��K���FN���PI}��^��)F�Uk��b�T�Xp�KB��6�j��:ڔ�������
(�����v��6T�Wꀳ[����%ݯ@�{JUq�g/�h�0�Z�f��͜:,O��tHW��O5[��*�H�� ��W⺈A�H���ږ��%��� ��u����]0���Ub�j�p��ߘ�U��>�����J��f)P$�or��v�-8PGӞ?�'�o�g�[�^if�e��{�:���]�ꒆ�}����<+���:�!�[0Օ(?+�o�U�+YɞHta�W]<��/����̓�_�[�����N�w�ܫ��� ���&�(x@���1���������+yv;޾�f&�RʈD�I��{Q����2�Ԗ�>���E/uq?��]+�����4n>#?1���BˋM��^a�G�� |�b֢��ӄ�E��|6S�m{��A�e?��9��M���ߜHlQr��gd��F�.d������$�r[v��?I/L���w��`��Vt�4V3��U1YMZ��$��y���uXP��М|7ѩ]˜�s&����A��%},����۳�����Da��]y��a��L��l6���W���t؝lxy�~���"���2MÒ��'�b�q�R��MgM���ZN��m}�����g+O#z��8��'jqg�C�>��WT�J��q�P	�����u��K�9YP��P4^��>�����`Ϋ�I>H�F��CS��G���`��oz���ܩ|^�q~�=����������<>Z
�]F���l9(p�K�8� �e4�Ѝ��d�W��(-�y�8\vP�bo�R���g�x8�\Ș���{����}�8��Fvѝ�GTɚyd5��T�U/�>!B��h�� �]�j!M���2�8�Q _F���ދx���O).���[�.F۷�'aT�I�� '����e��;"l����|�Y��T�	�oF^0{�1f���ok㘥�M�
�����~`Q�0VZ���Q�z�e2z1C�(V��[�N�[�L_U�v���g�'��Y�xͻ�EH������(;�����4 ��]o�Um�4n:E��0�Sd��=���/�<���Z�cr��=:��'��L�y���A���]ߢ��U���oߩxy��� z���[uOM�T}x��۱m6U��Ywn�����l@?���ϕ  �H��
����z��A��=��F�wB%�ډ��)a��Tɒ78ѻ�Q�@]�BzS�
,��8:l,\{�֦�k\	}�ԑ4��mVU��=�>M<[�a�GR�����*�����}TS%��V<}W�	����ހhݿ!�v/���ܤg�6������AT�Շ$��(��$ Rx�ՑeO|vAnqV��jy�.��p���������%��5�c�B�hdWB��w~���?�o�N�k2�m �0�=#����_�GXpn���V�_J���v��X��_�ͣl� �Xwެ<�tsV#�>��{���|���1ӝP�����/�|���D%O���(]��Iǃ�������ș����%
}b�o㘃ˋF��5���\�r�|C�Y=Z��_P_G.\Ƿ�ݰlٽ�(RD��5'x�C!�g�8���oΔ:$F}"q�#=w���0г��&nŠ�kz�gX7T�7��wIo��w�,���H���a�9:ḹ�_�U�S��PD/�0��0!���}[����/��J���_Y��Ҿ�?p�*��^��e���V��+����u�^��Mk������˖m,��<���$ �l�~��_��s�i���Ͼ�j���$��t��fa�/M��w��$�f.���Q�3T�-}��Yw1H�m5����Q�W,��0���welH�mx1� �v�l�����#/u����y^`�N��aޠ,!�s�P2\�r[nV�~���h���+���\�����[������-�v���й#��uoN�U���;>Z��]��`۴&�R�x��H�N#���d\��-؃eb�a -�5˽��	�q}�]T*M����B�Y�u��?�Q��Rk��ɶ�r������O#��BQ��<;���FÛG�æ�?ivԐu&3�6kSۄ�aI��:�_���u�|S�ѣ�{8r0��S#���K��T��/��u������g�7��8^)̳���Q7ʎ<���$��t$�~�g���I�D9Hͫ�NY�|.:+ɞ-Z3�\�����ٓ�y0HgZŔ߯�{tg|z��q1�>����}�eSf�ksAݹ!�d���!�v����:��B�O�:�o��_����@_��ng��4�^$�ɼ�m�}ܚ�7��E��>�֟�y���D��?�0����_Pw#�Z�m���;t�^���M�R��l��]V=[)?>GK�o�7�(��;�ː��E�?�'�`�yT��qo�'蚾ڀ[k<�8w��[{ uԀ�O]a'&e�5��j�� �*o���&遄�^����~z��p�D�/�9<Z?*2�֣i�7�L��&�\TH��C�����tyy�՗�]qqԀ(��
i �_o��'U��"J[.zyNȬ1>�LF�_<�`=�(����`�>QQ�3��&�ұ���_ԯ���]�)&�l�偼��ݴ������.��9p�s���%���qw��k #�WG�>M��Z�T~��w��z|.��Ȗ���c������tB�M��S6�)��b�'��������_�̩�9�xQ�{��b\����#�C7�+u|����l������x:���ܒ�[��SՓ��o�?QQz�oH��<r <S�`�ӡ�^W�~��;��1O��nUyyJ�ۡݠ�g%��ӯ^ࣉ���azYe���R�Bt�͢|Ie�ی��z� ���0 "Я��5�[�t��I%�J���'8�Xݓ�B0��{:|� ��W���n�>s��Ff���m�W�p�;�����[�E�na�tw�0H��t��HwK�tw��� ҈tJw�tw��C�Ψ{?�~��������+W��Z�Z8�~?݆ܲ�}u3N|�ޙI�P�N��-�|��'��pM�I�M��v�7�}oZ��ƴ��U�Rg7���$�&���ж�>�L7��-$��&�+<��w��'<�j"ˁ���%�ObH�#�1Om��Eڙ^�`��<�f��k��\��eX�ua�|�4N�=��xdh5Y�q��K�X	�ڏ��u>7���q?��^*+���8G�ڷD�G�?�.�Z��R��nRYq[�'��ds��/���1��^�)�����$$���~˩f�UɃ8Z��׬���/��L��M�����9����ͥ���Lm��.����R�oR� v#^kq��i�3D��s]	ڜ~>U�ַ���.P��\�5�i�1NX�e��cV�WO`/+��:=HE�X���e:�"��X\���x��f;���<�C�~���U���g���EgK�^5p��	b^z���G\��O�����=�3���D�C9^1��vo-�s���z*N��scv��JG���S�&V&�A�P�b̪4��o����@[v0�wg��U��w-r�.��[?n����l���OLW�>^I}|ĩ�D���YOD[dh���������#M�����4?�'��:���6���EÈ�s֟�FM��cu�zn�ɦ�ES����������?C���O+�Y ~����h]�@����>Թ�44�(Jޕ��d��}��K�)}y��
�K��xW��ɔ|����`6IBM��g���Xr���C[W��B���8 ��*��e�e����j�"�yp��?� 2�s���O�U�A�Yɬ��D!܋�-X;����~��[iX�X�I��(��ь���£s�t�S@�4�`f�G���;�?E������'^����>,�I��й&�;�������h����2g��w�a�aZ��}a�C��7B�������s#��[�G��*c�3�����)�;T` �M���ې�eY��z ��"��	r�T�m���ب�4|X��zF^*���$����~9��yRx���G�{hg��ш��OCVP�'z���U���T�������p|��j�s^�}��H�"M�&�"���a���QM����{�Oװ����?�#�0�oӯ�Vx�R�{}2(�J�F}��[(�ZqPb�,�i�2�VKN�}T&or/�^]"�He9Nh��`���LA�e-�����C�{&{r�o^�w�"�Y|l�`M/�!2�=��CB5|��b hټ|��ΪJq����Ϣ9:'�O���-�l�-�*ҹ��Mpm�Tj?h|�<����}��CKy^�L������Te��3���~�;��ʮ��d7-�䑵�T6�R�)��CgE%0Lg��=,kQ��2��?J1����n��CҔ��&�?)�i�Y�T��Hn���oE�&B�e�x�?��k�:���W��+phWP�''k��]���b�gw�a��?� RMǝ�lų�AS�H @;}��<��dm���r�,�8u7nՌ8�Aꂀ�>�7��? @�۬fP�훡���)�P�����X���gYQ*W�s���Y/�����9`��x����9],�p��~��E9ݠ�W!��hs�gJ��<�V�>v��&9��P���R��yBU-�߆F�+�3p��;<^v$�m����.`�ML`�-s��� �>�/������2��tI?57���|�pkS(�����T ;���Yc��z:S�9s4}j����hN�U��B�(�x�"Xe���|F�В����e�Lpw�Pi1�:��y���wo��B������k߽T��A��vdg;l~�l�d�h�߀՘�_ŀJ���ev���A�
Y��&L��4Dv�����W�d=Ӝ?�g��	��=|�I��{�ux��^�^��Y%� D����������|>��H��6B\�Bm�̾4���ī�*;��/1ǥL�1QThVy<
�|j���UD�(y� &�>@�ɗ�`̈́x�8�����G))/������ܸ &lEJEf�=�:��ӭ''�]�M`�����D�x|d˄�e��G�%Ϳ����z��K��T��ç�D��Z�k�Y��؛(�_D���x��\��d����\��oj��8�>���U5 �����]7�gl��¤;d�����|��22|~{��I�Mq��ag���U�7��r/�ڈδ��N��4<p�(;��K��{h���Dw$���s�7�6*��%�R74Tp��1>�i����X|�������O��P���y�1u
h�}\qYj��c$��K��8��+�f�C��1�&B���ʯ\e��{�V��g�d�{��Z͖Ƽ+�p5����<T��=��J�ʹ�L!|=� ���(*��N�o<rA�O�[汚W�}�;�w$W6}]����ص&�>��@bӧ��fy[�X|����F�>6\Ar�E	vځ	OɘX���'�模.�eSl1��|��W��ǲ�4�|+�7�K�n�\{K�%b�3۪���J}<�{w�C�.%��r?UDl��F1�M����a���R��ң{�6��f",���s��x������1Pa�ڱ3-�<�bk ��c��榷5G�;8m:���c9��զ{��V5H��\ѽ�����ܟ6q^��+�%��HGDj ݏӏ.��O�{[�ee"��)�N b-�0�����?,f�BG���b���q8DG�d�GK"��c ��	���~�e���J�*���q����;^�}2�2nI@@K'Ӎ�Z�@����֎��G�z:е@L�?�&4�y�u��;+��^�7��\wᱣ��h�}�!ea3�H>��z�GJd�)�1�!-�p�����(O� �W��?�Rq�+:͕���r�1�|?�X����4k��pd�fS��K��Dϝ��G����r)��MR̚�h�.6��<i����yI���w�0w��<��NӤ���G�|o���X���_�k�R]���B�d3����(����Yl�}]O%�sq��ꈜA�W����W *4�}��2`����H��;�S�9�gq�ҰY�d���[�l��فEoybK�-��!�}��
�sy�\.��<������!5��h�C��)�)���D`�i���?�#T$X� �U��E� |��髺���ڦ5G��+���e�V���2s4�n�V>5�	d�X`���z<?��y�k��s�6Rڽ�����ׅ�UWV��G}ET�w�� �����.f�'�+U��B��!���ҟ��P�+
�@��f����k��.��{/�T�PT�d�J��D̥���:��B@����/���@7�K�l�h�4��*�~���P���t{R�3���.���8��M�Ф�w���l'�oA�.�g@)q񃱕s�_ϳj?��hu��C���n$�x�h��fY�H���������ݿ�� ���e�c�Q�e���1�߉�p2#��������Yq�+i�K�Η_M��;H�
�
=5ݗ��]Zh���Z�
�&};�9�%���t�'�Z��Bͼ-��68�j�T��cˋ,T8k��Y<���y�T��E����ժ�d,;�q�a�@f1��*m[�?�4��g����܍u�Y��~���ƹ���<ö��&����юY���kmx�z�xAͤ{i�kd�%h>��s0`9J/�c�T�m�Y���(4렛.�(�kk~�+����T�I½���O���K��E�
���i{g���g=WUN�R������ @�ӽ�UL�����"��B�3Jud��orZ�J��[3.B����!L� 2PV�n�X��靅I�m�կy�zI�8��,
��m�f�hPh��*�2�Pj���>U�v{x�,_�ej���rG����]΁˛�}�E�#t�6�U�~��.?�H�T�*p��~B[��_��8�A�)<�311�=�T���g���w��A��ڵ�'t�eHs���b��b>�iSI��B����h�/=I�W޶�@B[�\��D�N��u�1��Pi�96�6T<����2��t�xu~�n`�Y��W�v�Dxk�8���W="$䴥Z�j��?���V�Y`��H`q���-�z��"wC�qIs1C�:<�Ы��B=�����g��
}-�ƨS�}]�R&a��qc�N�i 2�d�p���޿D���!ľ~c6D�"��Q���a޾M���V$i�m@��G8�RM�i�⏤K���Z ڳx��V-���=3�OJp'�|��g*&!)2���H[``�.
-�p�H�P�d��փ*��|��^��[�>AɮK'��ު���?��߁�L ��Q ���j˲�p�X.8���*`tٗV����;������ѹ_{a�A��ᑱ0�.�=?�����_ѭx���y<n��X'9�e��C��(�An�t��1�x�n���{i=� ��Q�"�+b 1U"N;-���S��@�����èK}�s���¬̉&qE�����s��{��geH���=�c��M4�?6F?,
��;1�8DV����Ψ�	9b�r�jU���z��Y�i[�&;�A�����{�"��č��ʯ�vD�2���zV�`D^�!b��pa ����l�zK��V�{�+ڣ��`#�8�j��u.�S�`Y�*�_:+���ٸ\-�x�L�Tv�=8)=st �P9��2ƖT~z�\^��G^?ك;DLQi(�[P{�R�����1j�Dj�.M0[��Y15-�_�|uW�b�|����Q�"��]���%7�z�H �rA��:�2{��E~e;�I:W^k@$�hGs"^ǿyX(�W�����r�&
����_ǣJ�[�`�P�7��c��ǐֲ2!��$�V��#�t�'6w�m[�d�my��ۆ��d�ښ���ӓ]̾�S��0T���s��Ҕ"�`l���9U$�O���)f�	�y�}��m�� �YD�Ym���v�s6��|�H�Fh��9.����\. ������w8?lg,j16�h`D�����Lj���`�*����0?b�G�A�⒡��a�Grn�ǣ���ܯ9�f��Ɉ*�SX�����_\�����0�%��D�4~|LC�_d�S�q�r�p�|��u���b:���K�swr�E=�r�
u�� �i�
�c:�ܟ�`��E�&V�4�BA���#)Ke�_�P�1�,�X�^�K ���/t\>M|�F!�ڜ��\�&V�MJ�Y�ɆwS����Q1�,)_�I���_F���v�hz@���w�$g+��rOI���
�y!�G7+��B̼׈�������b��J�gs�>L�Ö
���j}�����ӌ�C�Q�Y��f�	h�6�Ї���~��3}pZ��':�a723���e/@�j�����K-�5�/����6Ph�7n8�;����P}��Fɐ-~�"����z�K�7Gc
�3S�˰F6[�[\%���Γ����g6��Y�z�b~T�k)n�;|�6X{@6ŧ5á�8��1��#U��j�=��/��/����Z)Za����^pc��l�K�d�nP��*^U�R�&+f���Q��>v�#��M�QN��$��:�,�7��c�]N���p���[�-�0|P���/�ե?U���u)4U�'1��D�\��8\x-�]�@jd��@�X���[DNePy���N�~��*�{���	��껳�|w��sEGǿ&�ހi�H�,�{�+�ԋ�����)@H�UBҿe1٘w��퉞M!F�>b���Ȕ����י�%��gi]-Zt7���	>l��ډ�����x�k4}°��=	�.��-f���QE|N�����Г�����<_{���iN�BcZ�x6]+9[�XEH:��S�+�V,9�Ͼ8>�/�`���?��·z�<3L��@E�R�P�'��J�� ^��H�E�	p�t�} �.�0�.J�Y0�(%f�$����E��ώ[�u�s�X��\�Z�+#�
ط	�[|��7ATL���(!��U�'S�t%�y�x�������IK���?�lP��{:����d4b�ĸ���Q-�����B ���s)4>�6}H
�{�h����h��<�}�	�?lv���)���T���O�H�`�|!&�D���TDOur�~U�?N�����'��D\��˦�� ��������L��P.6}8�P�>�~�q����z�����)߅$�*��q��I�N���/��v�FQ5��%�ptm�M;�UFX/	_(�N��D�MzD�cq�0�~���3�⿮��/����ٙ%{��6���M�DaF�h�>Q���1�g��R�F�K�%1ʞ6oxMe��][���}h�R=R��c>|1�"Gb�?[Uuy9٦ut;��8	�~��;�p�<(R$a��m�|�M��<����:-/�ť<B������5!Hݼ�s�n���Ѻ.*�g��e��U�� ��7� ڝ��\<���~w��Ϳ�T�ȗ��KKFdI�,��~8r����\S�Ju��0�b'+� Sx�/��nǷ�k��%����(\4s7`B����,vv��+D`v�v왨<Y���ݭ!E©M
w��o�b܂i~kkem*�'3zi,VQ'&��GjU�W���������9�1����O�,	��﨨(8�m<}�-�$�7�p��7QY_��ǿ�aM��rPB��Y�`�T�:�j��f���翚��a�j�T�vz��3�_�ݿ��!��v+���C�PZ���q�A���b>Dc�X�N�Y�������10��Y�p�~�$y)QQx���i{H�ײ;m��zgm}h�r<��<�ṡIZǩ�Ts����1��#"�f�* �b~�|����[J?�a�X�E����
1m�ЅDv���C��ߐ,�,�`ː��Z�8r�2�g>�V.*gp�$������Q��a`^F[��K�M�'��,?���oM �dO�l�N�� x���?j�'��PJ��TvC���P�~)3�g��	`~:����m�0`�zT���e=ܦ^����-fn���%8�����`�-�ղ�0!9@�{������	*�6�(t���ّxV�?��n����9�,���՚>7`ޥ�u�=4�v�-�}�0Lt��S��&9��������s�����^X#�~�.B�u�(\�B����|�Y"�&D-w���KIT�fr��?W��T�m	�6+�/�йB���wt��Ǩ���ZZl[l��D*�-�{*��T�:�%�P�~q��Ck+�P��t��B��~Wf}V�������q�\�bo?~�W������mN�4��0'X���M ���	4�~�!`��#�9��Lv$E>cFgt�B\��4�5�K^u|IL7K��/��*W���P��uI�Y��ϫEкYE\kC���1<d,S�&a���R���G���fF�� r�_!�k&7��N�]���L3����5�heϱ������[ ���p��s������g-��!t�J�pȰLW���}/J�dŽ�����ȸ�:>]������ ����L݇M��/�+���߻9U֭m�q��s�<�Ӏ/��T�`���P�{��b(Q	a�a��P �"�,n���������I��ɛ��y��k�TZ�!��رtjWP��cs���g���"�M{R���֨RHcF�^/�J7��F�Q�����3��p@���O"� 1<��]D/�
�黥T$��O��4�~b�N�i	����?�.>�-�q��������ƨ1�Ɵ��Ь�n�uK�f �#��^��6 j���T.7��[y��ϔ�2�����V/ᘬz�?�h-3y��aj"��~g  ������r�Nrk�N_�B<MıDͶO`����(x^�6��xg༷���K	�8���[U�TV�!0��_�]�*����<݀�w�*GVVDJ�8:o�4���{0� �p�oM�t�w��Vk����+B`U��͙��eGg��{���Mr�`�8�l$�p'7k��if��c'e�����'��u�E�24*�����XJ|"�?`�AIR�;�<�ո����Y���>|/�(\lA����{�E�z���ݡwi���i�5QX�\�~Eџ�U�J	�����A�_d"t�D��A�Ⱦ6e��rC���s���ݮ
P�c���`���zn�F�oX�.�}���mJ2^�� ���.�cG��H���0�ۖ���Ì$�Āl�Կ���� .�~���d����u-�5��'��N[�
i0OF�N]�2�ǉ7\�b���M3������j��/�?�ÌB�G�Ş!W䮬����������7�c��i���#�!,�Ǆ.vEƂ�@;��`����!�6�����tl�2��@���K�Ԃ�!��5�-���(	)YWH��i3�iNFKo���~	�cߝ/\����"�:2����{^���®@�(�mM���|��_n�7:��K���dY )�i!|{��s���(u���V\i�T��?�4�Λo��:5����AU�02d��r���IOy����Sk3T�\���<9��B��[.Z�����z�� �tK2���N��.�ƱW�o�.�b��������Nʔ;�E#G�J�I�����C�;w:_O�l=��8���9��0�x��={I2��a��9�+ͨ2;����������#�K�Ӡ�Ҍ�O��I^���a��~F���Y�A�BOAό�2��c�e�o[+�����[�u=��!Ճ�"0�eń9#1������ DܣD�*^z���;����*~|�_g��(;$�W����KE��hSi��{Dy��*z��G�-���-��mЮ-�AwS0�#V8�����~������Y
��<9,����_z���un�K�bz��49犍��;����g��G"?_bX��0M���2��J��ҟp:��H�숄j"!FUA��7Κ��Oc��;��t1�&t�|��/o�ɡ10VT6�����䟍���.k&v��n;9�vTu�(�u,��T�'����O�������������`��)|���Mǣ�*��'����b��:���X(�؀���|߹kŞOn���W���I!3t�����qԦ�}�����q�����=N_�l���2Fv󜛙��+�U���G��΁�
�ͧ@�	�/���[����3d�)s �e�i�T=�S�"]���&�!��w��y���GdN�^�4pلO�Q?�Q8�N<�/�P�"��ήm�7���P5pj��_Н�/�M��mP;�����N\���XPi1��Z�<��b�.?x�}	�ED�,}x��M91)cyT�~�Dlӣ`�e��4A�*�6c$s\��a^���[� ��}K��Z��M�|������t|	�
��'���KW��6�p�=\l���1.H�do�������YU�3_W�<L�a�'���������ec��v�;([�sW�zP�����(TP�n)u��+��M�o���A,��"��V"����j�MG����Qv[�q�.��[�Ǯ�w�H�e|4�H.v�H�<�t����)!'J}P;�we�Ok�yqle�5[`�z�\�J�{ �SU	.,�[_�,��tu�^3��	`URԽ6q����q�x��M��ePN$I[������QeK���4���yU��^j��y�sQ�QV@�B����mc8ס�R���⋦��E������09�T�qb�GC��/�{A�e�ZTG��<\�;�G��$����X��;w�LP�9�<�:?S��W��Ҍ�G�"/���7��sv�3{�[O[
��5��e�]��|<�
�z�,f�{�K�}s��๱���GmsP]�s���|�+���C���%�������Y�N	���o����+��t��O�|p��UI<DL�82B�qpgx�,�ȕT��~ш�GL���ȕ�xw��?� ��}��Ω	��/^��Η\lD-�Єn�O��MCt؁���.|�3��pS�	��4�sw�W����/W$3]9����Gi()1�8<D4�S.��� (��ź<I}���Q�c����6��ϔ�-�3�աZ����< |�X���%�DMW��X8�����}d�LYK��x_�w!B��)���I�ɭO���`�q%�,�����kLSh8VDc�xB������@�����7�\������k\D��8?$*V����[�'
�@�S�"�Ĭ3���_~���h[&�{�=v=�4c�S����U�h̉�q�G������K�Z�"_�
7;jN�MS��ޮ)s�`��m����͌��nx�?=M�����	��	��X��1ѢP$���'d� �O�=�c�b���o����^6Ζ.ΐ�\��k׺^H)Y0�����d|oP�#B�'�Oz����s�����qE�����zd��F��av\sS������ʅG�񛩃I4Z歒ꂼ�g+�ĭi��4R��wd��Me}������`��*�2�G���)P>�_ ����AR��bf߿X�k|�5o�.JME��r�^4���J�Үt�N:o=�7���Z-M�.�|md>^[�,^�!��{G�Ęg��JfUR��Z5��gK�c5o{�T��W�-tn�A�����h�c�3���%[h�',ȸ~d��� P�;uF��F�=�%��u(�'�.#�r�2��w�aw#��4���|����� f�Ry�D�_/ز+�Qy��p�H`9�5��G��Ŧ� ��*oi4j~\q��DA󢡚�!+�o���	�
�7�"�ǣ����tT�|gC.A?x?�<�f'��S��� ks��	ThZ����-"����`�ɏ�s$�)ᆈ+�xD�R_��c�'�ac��de�i��%�D{<
l������n�/�z��%3�V�C!
��v.�0����
n��~J�ː����k��75��D��]F����c�d>1���[�=\��&?8�`��$���v�-FD߇J�ө��8�;��ŭ��RW$�NZT�w�wY����>��r#�e#�銨����^�m���{>J`�LW7>�^�꽦���!����G05`�BJ���v���	M����p��J'����G3�ꗊ/&���uC��QgT\|���1��+�L!�3�������p��gޛW��V�j�t�m����-by�����5o�y�ޗ�>;�N#���?�G�cۙ��P72��ȶ�r}�P�s�N��~Jߓ�VX��"e�#�渋�������#*��Am��=��(���Ȋ�TW�i�o�l�Wx����m�$�V�+��*$h��wML9�ͅ�9�����^J�xe��I{�!Eɺ��W�[�X���JEH����'�,V�G���
��I52�@)�Z743�Ϯ4%�#�7���>?�d|u����d)�P�'��8��Jȑ��h���.�� �#��dS㲯�KU����'��u�	����k���w܅�����[(���27]9��;�ON����Q����w�p��"����p"�Q6i
=([V�i�>5��߷Nʅ���ulë�d_�$�t�q�@`��v׿�W5U������d0򺅸B���f'D}i(���K��� *>l7[��P�Dş��cŔ���6D{�`����J��w7��Q
��HVa<v��|���b���"*(oh���*->��PQ��>O���$�%Y]yF����%�[��$۲��N���/U��|���y�����UMBE��ߙ���I5��B}�M�Kkx��Y�(��n�P\{T<�O��C�Q��ˬ@9&i���K�g��(�;�g��E���=��5�J�wg&�G}CT{�xpL"�$��֏E��
i�߱��C������4Ͱ7����R��-_[��T�������Y�Jn�"BC��#F&j���*Jz��R�l��� 9Zz�ν3����h�EP���K�W��y��2(�i�����^����+M"cs��_6�X��N��fΠ�*i3J�'�!0=�Mvn�ѷ���rC�s��}E���2+F���?g���O��9�%�^���D#�ɬTCLuj��N�������6���$7"$VB��~΍�[Q����7��A������?�U�8�2��X
�:�I�&4�z��#@�����J'uV������p2O�
�?M�Z�~��0� ;���盀K�!��*��e�,UXx�2y��~��=	_k��@��*��{G�.�@#1���@Ʉ^=�6&�^l^�k���j;S��<�,l�����|����f
����Kmͧ���xo���l-����r�
�*� 1֑�M��V&�F��{��`~��)b�-���2(l���I����&3�Ͷ$����sn
�K��|�B(w���0p}æ�D�/�JƆ2�Ӯ*vq�k��n#���͹Kx	׆��Ƒ՚��B�"�%�i�2��4W��~g,P�6��jWV	傮t!\��К2U�jc44�~FN�vyחq�O��b#.�gC���s����
���%���8��W�0`�?gD�Ikn����ce��ɐ��$����(�,>����b�/���>e�_M��^$} ?�T�Ly�OϢ��ˮs]��"ׅwdYRҒ.�	Am����:��%F0O������Wɍ��S��j�k:<X��ώx�
q伞��[���0�v	_H�������{�]�x���5��K2��ſ*���:���&f��x�����η�\�f��R�?�_m[�໽��|7�����K��&�������H1��W-��}h���&�����~7���L����VE��l�	�Gr�>�6�dFd�Zrpd{:��\5Ip$-F]���xdl��g�=�Ͽ�
��K��$�g0�d'7�k�訴����O7M�g/	mzK�Ζ>�B�{[�Q��wu�"y��R��8U�4��>�6� 暈 �L^�����5���}_��uA�L�S��o��ؽ���6�+����|$ү�1���%cr��ybϕH;s��T��OnOz��+�H|�zr2��7nt����'����
�L�ڃ�1�T}�W�r2���k�c��=����m�T�@��6�\V�N!a=Kdg#/_�M�M�!@�v�IL�N���O��h�>�������\�a/�h�����OR$�e���y�:%���a
�{K��U�gɓcAZ�ڽ.j���+���c��}�G�� ���~�bǑ����j�)G돋Rn}D6}^���d.�#>@��&L}'�.'���	��ᦍNF�Z�������ɩ�Uð�X��<[��MMI1�2S���z���-KVa۝��8{}Ø<������Z�ᥣ��bh��!��C�*e���'���e�� �o?�Vi~["8��m�>�)��}?U|KP��v�⁠@�N�8 3{�.�Ol��=�ׅ�l��%���[�N�ZX,X����cڗ��+�}#�����>|}��F
>��k���8�u�"� �S�YD�!���}�Au8�P��w�X��C9�p*�Lq�f�=[���K0�7+w�Q�B����J�1���=��*%�o�����y� ^w${mW�޿5c_�n��/Z�󲛠�yl7[����w~�RҜ�CT���N7A�X7A�Q�V�_|��ն���?rp��i:|�ЭR�B�`�`�̶M��T��@f8�/��/�>w_NjP������|��0�fQU�ǁ�L�nYL��m�M�yU������d�YF��/Ԟ?4�������5��]݇G�������-
���2��s�Ta�{�>23����;�T�F���]|���1�]���~��UN'�i�{��I�	�@�}�r���!u�Mad�V���Ϟ2�T�Ω�Xe�z5u�ic.�j_�l����x��i�D�e��#�t���h��G��N�(艀U��;�T4
BW���J��]�mb��Ø}6�|$���/���	7`�2j��#�cו�+a;?͵0�<��6�d�?�/[�X7x�h��0������?C8ju	����$��]<B�a�
Rl:�dGJ���*#u�8PU��>���+�^�@Cf������^"7&�2������*6��2-�@�V�9�����[<�r�롎�����&�)s_��������"3��S��ڐ�Lȧ99uO����Be�Ҽ'M�C>��3k��ZՏ0-f6��0�MJ��5ri	�MGD�O�|f삏�]QX��|���&�K��	&r~o� -�u )��.z�%T��4����B�� �������X�["�<�Y�w�H>D2O�353i��8N��+pd4��x�$�<�d�XI7�6ʄ��J^�0f�|�3I��l��hH�
�]�j��j�\cGj��+^C�"���C,��D��\���;��#�����={�/6/��.<�)�!��+��{YS���,d��j����p�Ǿ�v�|�{�aB�K�P�ă��������J�dYŗ�ں>�䨼�M�H�I.�l�œ0�ny�D1�1;{���N�|�j%�v�_�����5n�C�#!�ϴ�>2A����@*�$�*)1�u��kK�߇)�G�vv"Y�l���y�k���Pfr<�E�B�N���l��#�Bɹw�z�͢��J��g+|�^�hb%�IC�O�?���ɴ���򊪫��C�2`>>ǬÎl�䮪_b����R
a�D@U#X�̫����E>����	����H﭅K��1���6�~��mT���:�H��0�Gb���v3���B�9KDv�^i��P�/S�Y6�5�W$�A[+v~��ק�o�ڏ�%}���B�C���WJd�U^cDE���~fȅex�i����,}-Q�r�a�X�Bwt+!���P0'����}����b/گ;@ˈ��d������hķ����iYk�ƽ$���Op�"2��eO��¥b��5�u�8�L\W3=%���A.����'y����|�B��Ԭ"�b��q�R�B�Y��t�'���R>L�mTRc�w%�(X��s�Y��������1���;�CD���b��+_�>��L��u*ôpщ�^V>���M��D�BZ���#��Az`D�OG��¤P-�!��;����'���>�ݢ��3�;]qF�B�R�z��9R�.I�vS�'Qވ,@2���y�$O�p抐����@t*!ݐDQ�]]�(?W�1�5�b�]A3]_����7w���*[���HX��:jŘ�A�لa�k�7�!PO�~��$�����Y ����i����pC_.�K��WD��%/D��gXUrj�����x;R2�Y$ �ﺝ�Msw�99��/3Ϋ�c�ޭ��+b�5 �9�;��w���#}>9�+��c{�m%�6�5ܠ~�-�����\V��8��	8���R����{'�U�q�	��d{��*!�L�{82l&H�~�o��L���Oǧt�IC�L�)b���8�KII�P�B#�:�����3R��d�w��6ݏ6�yϼ'�'w��o�W�Lʥքx��t�s��T�1ȷ1�͡f�Ĵz�uS��F���g�	���on�Q��sU	/P���9��~��޺�p<x,j��Ǔ&�WaK����7(�sW��|R������|��뫝Mԩ<��M�	0��^����K��s�|��.T��:�)�'����UM5jl|n�V����Fv��3jn|jn�h��?��[T�Vt1�B  ������A2��\����m=�6{���+��-�������A`f�u�.�B� �����1�V��&�B��� ������P�<Ӿ���@���0ŭ�LNg,��W��,Z߈�xlf�?^�����Ʃ�]�'3��uW��=��c&��*rK�|��Q!E��F��\�s��k�i���.��L�.���2O.������I�J�KLU��I��Rx�g��/;<(�4��^{�W?5�x}���ב����|�����u��h�=/�~ga��O�4V��	��En��)��a/ctړ���5�	��F<�~d��<{Z_�|%�B�H%�!��Mu�D�<M���C8���S�=���Ҋ�S��)����"A �\�J���P����'y�Q������mo�
��T�8^���ؼٛ%�s���������l�CQL�_�0&wb̦_�3���"������g��{<D��͒������2��5^�5��
e�Ya#�Kh����b(nK�>���2�UiA\|�Ӌf�ښ������9�a�O�]�@�����sf0w��Av�f�f�2�&���D%ZvC�D��K8B�����@3�Euj�Q&����V�jZ�=`ro�d���I� O�(��#�'�B������Z¢�c��p/DV#��|��`	��Gq�v	b!gp��}��G�ݖe�	?��4���]�0ރb[7�|�tE�><��ԏ���ƙ�pw_�V4�eɃ�V|ϞK�'�+���x��b<?~l�ޢ�@�Ψ!U0Y�^o:YY\>���%�Ŋ��1Ҿ�i���/���o��~?j��R!o����q>�x_����3��R��#��U���! ������e5�S�̓������(r�hN6�n��O(���ߓ7��~'�����,���W0ͦ_+ ���,oŽ^�F��b6+�"A9��7�w�f��^�E_�_����^
�ˡ%VG�R��4���ۮk�/Ь8ڄ�?C��ib��u�-��O�%�v5�F��l>U������a���=�ۉh��n�{���"�����1z56o��]��G�mF�څs�Xm+$��,=(MlK~.I���Cg}�:ӿ6� y�ʏow{��fZ��o��v�f
�: ;m�׃�?\�uX���>LwH7l$%�� -HwKw�&D��CA��ERJ��;7�oo���y߿�.�>{�̬��}Ϭ�t�����*$�碌ꌪW�ٿ]�� dY��8ޗ
�Q��޶V:j��<�4sz괞�{�����AE��d̫Ʌz��볰�*,h��� j�ĥ}b[�AŰ�(���Iw{�!�Q��"x���Y�!��X&�g�o�|��X�I�~cXr�ﱞJ�V�p�s��v��hˠge)�:g�`�C$4��oX�����6��^Η�,V�'�4qCrO��V��,{W�5���-_
W���`}n2�&����bݑg��n-�?|����1�"`?F��!� ���]O����L���hh��HR��s2�	���m���M)ɌV�Xߔ:�lvT��Y��O��5߻#B�SL|�)x�BC�'W�%mq�����	���I��{���y�lo��Z�:\�i�V~�}��&�6�ٿҞ���"��b�̙X��7B�:@@��3��֒O�����|��p�(��*�?��P��5�-�Q9?�A���B��	��U�r�v�~5��n�j8��>OP��XNl���ð�꩜���"���5���ĄZ�cY:7*��3W�+��\� 8Xb�=� {H
�����!V7iC�J׿�,�Xƻ�MFBΆ�5-`2����0���x�=s��Һ�v�Tv�c���|�2�x8|�>�*���c8/4�9�Q�����S���+�=o�q N�}F�2,*JA'(�{���^Ǆ�1>�'9�?&L �Ԣx�+��[o\��g����'�Q��=c�F�f��X��ڤ���1��8J�)�W��{�D:k��	LQ��M�*ۺ@�l�?����|>ȢNu��c�I,���YÑɡ�B�o���_"��0�����͓��i���b^��U�o.�G���1�J����dLG5aV�H!3r�s�����)�d��;?��~2P�x����49 ��ߍ(��L:�� A����(2 $N��n�,)鞀a�_��<�r�c�bt�̭��F�s�:���Rn֤K>��;;G��+�oë�����u��҇�s����}1��^1E�HKn�z� ��c��儙0��)o�DS��o�ہka�wNc��s����
z{eN���@�B���n�`�`�@�]#;iw�cI�('Xr���L�L82����(�!]�I�jC��qw�3<��0+��u,/=��5���aHu�*ŉ�5J��f!]�@�|�]�F��s��7��0�3>~d�/1�*H�_|~�Z�/�OI�f��@��)V}�7�}��{�!*�89��kMݦ�HU� S�����>����������G����$M�$�����ݼW�Bs�cb�D�÷u���GK���A�_�9�]Hԯ����~��@9�G�(�l�I�:ڳ�aY��:�Tg�s&5W�Ӗ��ށ�T��uq�%AВ�Il�a��DP������na:��O�/f
��'���I&�S��Z"�t���4��u6>k`ly7�����1�����g�S��,�L�3��<�sO�q�P1c�"em�`f��}�ƭZi�8�˚�;0{o�ʎW���@���f4�[D���-���X�ߏ���cC�2,��3�.��f�/,����:��d�ܕ���-c��3Y{�fu1b,��U�"v% ^ށ���z筪�{�*\	�+� APf6<���\^1L����I���Ā�Q� U��N����4S�T��J�@�p�6?��~�	��|1U� �[�l������a���ӽ���ղ�<�+R���q�������O�߫!�'L�F'J�7~����.�f��������U�Lss��������IkDr�����tܓO�(L�G��
� g*��cx��1GR��ݦt`'�Ti�G�(ɯ���ސPe���v��97r8$ X�|�����z��@�������>rMy�2˔qɝ����o��mJ��u&�˄��*q�3%i��|��`���\�a+���4= C��*��b���؋�q[�74Hs;!�x�L��
bq
���ʯ�=�v�KJ36`>����a�h�
���ͦ��������L�0`'�W23�2�����D�{-�?Ѩ�(l�A��A/�_�RV82���D24�d�cm��T��z)�`�oS:}f�GV��)7Ⱥ�}��$獰����ѫ����)g�u��]֠��P��6|�$���Q�)hx��B����5b��k�N�(����~k���������dv�B�"�d1�:�6;�G�?~�aKNʘ_�(E�6cTs7ꖹ�^R-��� ��Ǌ���p-�ؔ�u
��p�\� ���*F��M�ݙv ���������R�D�֫�_�@���Ƈ$-������-u�/L)��B텢�c'_��U�ō~u�����)E? A��7
��>�Mk����$8�-�J��U�̳��W27�2WY��׻ߚ��$��t��1%&��4!��^�ߛ�����)_!_Ko�C�졵�ڨQ&�:��w��KKW��S�KL�ňJL�@�~��ǉ��FU���c��qe(�>�����Т��f���߳Ŵ7��N�&)���+q]�sBi���/L`��>�o�b��&��Q�o>n�� ����I�*+���k��#d���еf��⹇��(��/: ����� ��ǩ ��濕d�<�.e,Zc�|�}o
�h|���AA���:�eMo��j�R?9�L����iO?��*u�UV?���$�{͙]l�����V./�3"�tGFxå8,2u<n�x�]��P�Dw��Q�*q��c��LC�-A�D�1 B�,'�R4��˜6�N&����bֆ�E+��^D�`���S���p�3���рK�s�$GϿ�-q��<⣌(�ሂ��'���Ih-f�n�LP ���>��O�$�Û��̺�٠����;r�q��5���f#��$�hA�.���j��Y��ƻ�L�T&���w���]-W�"zJe-�gc�y�|��9&d�0�U�c��lG^�{8Δ�5˲�LG�:�m7���"pl>������P�AV��?ї�����m�|�h���A_F#�R#�dR1|���=&��W}���N�	d8��-��0h���;�b��j^R+tJ�o���y�ǽ�4���������]���q�ǚ�O�>:^\Z�VK˿Q� ���\(�^�2S�]:� �G���po@�(�΀R�W���m��Q�f-�9���hg�]�w�@��Ɣ}'������=���*Z>3n��O��B�]�Opu#�����]*�r��y�A���~i>�$@�n�&�*0�}�Ӕ=�Im��uJ�fd
�!���B;R�@3_/�3��}��
hlr&�>���5�X���I�37�?o;ft�ސ-	���7�9^�=�C�J8զ�|$��$LU�kCx��X(��6k���G>�o]F�:����"���p�%�ʷY�;�P>�� k�Q�
]+�7/_���n,)m��Z8��Ij�ɠ�v��=yfV��~>� �E-�X닽���=OK�f�65�&{J�rW�r�WN���L���i�aS���˴����*�ƻ;.\Q�46yO�#�d�O6�T���vή������G�$hU��c�T�G[}���#fx+� �w4I�H'��I.ʉ�߽\<�%�Ib��ǒ��}P��/L�������dF��_�!�a�8]����7��ѥ�!��l7aô�کG�
Nv�������<::���|W�#c���c���b�TG$KA�*�@s��7	UH�Y!(g�)�L��<:{�3t�-�F�S m�@���C)]f4�c����\�P���/���z�HC"�r1�
Ca�e�WM��!\�3������<�Ռ}D�m�/u�(Q`�O��Ma��ƨr�Q0�25���iG�m.z���q�TG��Ѡ����_�Bk�u_�. TlQŧ�"<+�8�^=)ԁ��SO�2ٗL
V�p�^!�R/��޲yp�{����j������9z�e�]|����)��~f:"Sz�PŁ�egZv~]=֍�Z/����n����������ѽ�^'�����AWv�w���]M�s����G(��K��3��=\�B?�g���t=��`�E^����,��C��))l��_yo�4"'���C�l��R�W�
��ux-Um��g�y��0�g���!�oLj��ĸ��-)M������&�F)��O֟��?��w!�硹�Vv����-��	@�c����,���T�f�։t@.�}c���}J�=��xy'
���Q'�ֆ��o����gh����͌N+���u;a����p�7��,=������N�$�����[m�rAhy�&�|���=�e����,a��zh�>$�٦��h��C�&B�ʿ�w\�h��3XzBJ�(��Y3����`����	nt����f�=� x��V������f�73��+J}u��<�H�M������Z7��2J��L&H�î
�Q���~eQ�ԭV�Ё&�k�"'�yn���zH�~������Y-��_�EAi�D6ٞ7���ڙ���̾���;E�>�x����ɯ�g�U��Qzܐ����$<|���������E�՘�O��[;ش^ax��s���ޒ��s�q?}.^5B�UǼіf��Er�=A�S���M+��ttg����%��ʨlx��R1��[e��%���W�Jsf��XW�~&4s�Yc`�Ǭ�"�ϴI>�Xݘ�r*�x�6���`y�S�M�s\L�U��׀ܶk�{�D�u7g(7���pk��3|�xow���D�g���c�$F8�QJ.$�����g���lo�f����N\�Ƞ�1��^��L)�g+�y���(������S�vG��d�u�A��ʉK�o=Z�Q�A`r��d8�C.��l_��OF�� ��I+5���BmPF5�hsV�ݓŌ�/�؇$"�j�ֹ�����cuaǤ���)<���x\����?g#:�-�Y:W�2�o+��%������=P%\}?qI�~���}�.t}�>��GF�16�6�͆��7R �fJ�d�|�4r.P���������8-���h�I�p/���ƈ�u
KA�H4�d*!�=�#��~�@4����s=TN��1�_y��Zh	��@��?fVŋ��H�p�ZV_��z]6(�z����K~��Æyrr/8V9�sΪ�Q�����*�H��I�'d�l<����b+�P�� `	a�����_�W�\9�Zim�E��;Σ���|���-�x�N��ץ�Hz���c~�C"r��m��|�K� �M;����n�ߴ�S�^`�Eo'���d:W�l��D�:�-��ܮ5���77̿�q=�t�:yHSߨ}B��|�f��K������a��ϊ��fj���>��5��'�#�	��Wd-}�����В�#a���6��m2��-v�XR��������A�qv�S�M��-�_6&�B�CEmTq{�@'o82��k]L�`�T\���AN��^�0IDL~=B
���=�����cp��tml�l�)��xG�ng�"_�* �>q^'�`��G亻��t��1��~������+ p
7�o@�)���(��.�[H�* �Ң8��QT�z��.��Ml"!�^�&Cw�5�y���=�]�}�w�EV�_(���TR�/������u!;pH�:�y�����5"?Mn��֡u�a!���grH��p$+ j�U���[�e�}�A����̎�~_�$�W��uj
�r�A��u$ ���z��^~z�3��9��<n��:��
�d ���Z�y��6	�q!&�����w�m�/�6��#z(Y�Bz#�F��;��TlEeڨ≣X��O�ވ-�ݮ����zs��T�3�'�M\:���>D���~d���BZ���m��5~��fG�F��&�T�ݢ�Ƣ�W&7���scK�X��H<W�=��^BO�mӼ-y��ш�C�x'���w�K��iϔ��Ad��[�a]^C�n_��b2�VT��"���ӿ2@ ����}��s~R�9ș�|d�w��_�������K-�Q%b'l2[&4�&"�׷��9�)�5�y=�C���֡�(���&T��o� �Z�]z�;�l�#�.���0TMk!���	���g�a�YwK��%�NT��!���l���2w\gu���s6<�9w�w���ȗ�����N0�m"tQ<_���wg0�!F�[Eԋ�㒝�9���M�`�l�� �{�Ý-�#�U�ٴ���:����!�{+l�-J���;e�؇|/��`��?��(B�c~	(���v��ĭ��~�:�~�h@��Hh/4jD��*Ѳ�^����&�L���������È:BT����p��~v�p��,�#&���%������@!Ɠ��!R~���46��o���q��~�8�!���Qg�x��{��z�M���������'%c��8!��ДyY	o�O�>��i�9P��� D��VT��_��-=�s���u�#�NXj/(�H�q�7z@�_a�N�R(�B�%9P�6�l/7��[�yX�x�cS"!8�w��d��SI�vqaM��Ҫ=u����i2Q��a�:���3냟����x&TG�����2�Ԫ�|N�D�Z���l�"s���
�x��yT>�)(�鲓u��M�B�V��򮡼eW����j����K$����t
?E|��D��b�����n�4xrWf�բ�|��$K"�V��Yɷ�q�y����+�?�vx���9n��w�?E�G��פaH�@�*Xq�N�!R�2t�~�	a��0�3؃W�OD?̡�N]5����,����=��Ii��Tg��%޻�nr×'v � ��?���[�%�h~��b��:�̈́��p�8��<����o�A��_�&���JS�Ĥ�St|}�?�����trjN�ٴ�=6�]���?ͽ�1��(���j������m��~X!����j�,��Q��f�����^���?���\���	��M�1�
Kc?_���*�����U��@+���^�E���c��܏��2���l���1ކA�ͱk�u���fKBFd��V+��@䒲H�P��Q���= ���Gk��ZWլ�Y���@�C�D�w|)&��9$#6����tD��	�(���-n�^ǹ�7Gw��ޮ͓$�[�7�f��4E���ï1L�s�#b��,7Oi�[�Q�O�BX#��
�����_�S�;(��#aMr�"�0(��-n6i�z��� Q j.�r��Lwj���θ�2���U>�zd���Yj�����4�Υ*r�U%Z�'5����Ip,0�y�����4�aƊ*�N�Qʥ����kR"h� ^@ӳ&�,�5�cb�jJ��	�*\,S���i"�0�Xh������๊��|�_�]�Q%EeZ֞+��T��.Xr�_�e�5���[�kl����}��v��v��N���#����Pd��>��B	wq��6Uko��`�(�R�"�F�s]�dB��b+��CYn @�Z̾ ����j�-�Y�3�q�u��ӏ�/�QL���V�������j�;���YM���?K����Ď̃cŌ�V��� H�%�2��`�s�{�~������vm1	��&���AD�)2sw���~���r�-�kג��5#z��0��Bi̹�X;�)�<�t���⺅,�8�~+P����uKz�	���C�@���1� �Ū6'3)�.��K��=��d�b�"z��*h���G8껅�t��_����p��I�;�
�m�Q��~�ؾ������P^�q�}���a��'�$��G,��C��o�)�p�b�3�H��w�ߥ�y�E��G��o ;�K���p�!~$�_-'�F�%��?E��q�HV3��@OC� �wLy=��@�E�����Y�-v�.��{F�N ���k`J�����O�����Wt�f���TT�&��c�� ����8����hM7Ml̑?D͈<���eȀ��+.�����8pj��E c��X�_�K#�<>�~Lh햄�X~e��(�:��@���7H�tNu�_wA�+רy�:�A��@�v�35W�{�[�0���	܏���$�ȌI��A�ۮU�o?��0~Xwj(�τL~w����b��<��t��ޟX,h)-��Off�F��JGF�^D�l�hܮ 3j}WU�9k�b�h�1�(��4���E�b$ͳ��<�](u�T��a��so��5��!���0�q�+�B�@8��D����Ҟ+6��S�J���$eQ\��6E�=�j�QF��<�@xm��UE��ya4H��4R�=��8��=�|� ��W��zM�7F���Sɶ�ӥ��e]��+N����^h�r��������._�WD8�K�T�5W��PA��u��������W⭨��[x8��W�,^���A�@(,�q
���-o������0�dF��/�{jϭ�e[�r�nvЗq�z���l��<-���};��i����XX �Ѓ��(^7Y߿�}�����<fҨL��$[]��b�#��q����&j3��G "5�r�B�u鬆Y�*B�}�ԵbB��-Zbb��Q�kcjN����B�����Q�q�!�9�(�jh�23:��h�+m��Q��si]���i+��c��4:��=�;8�V�[Q����/�U����4��7||�����2��-��F��Da:�����Z�N�a}W�ٻ�h5R`o.;�?t�j���ëҫ!8II?[Z��)�����������]%�ޜZ�^K�7���YY���{vÅ�.�㛏Wf���ABc>�v|�F�wr$��0��5����1'�b8��b��nN��,�q�hR�� aG�򬊧ȴ�P?Y��Z�@�� 1��]{_��� AE�z�>�n�&��/#w�";�����i�����L�k��<���4xx�v
R�#Q�z��*��(��ƍ��X^�%Sd�6���-�4+/8xǽa���{_`��t�}N��]^{h����?}�t/S>ƾ4k\���w���3���>�g&��| e~2�n��z�ɠ��B�M�J9{OW�&0S1�f�C������,vŸ2X�C���'
ے	�;�.t���s0�2p�X��|V���ۇ����Q�PU���HG ���A��^4�P�����k:���ܚ�L�,~����m��v����1 �L�iє�cP��R2L_�%�T<0���2�']��l�YJ��op�6>���eS^�vm\}�T���3��y�m^a�n&�Rp�@w��{��^1�V��(���fM&�wi�WS���qʳxcfa��[G�?�E��/�6��L���i'�G�Ⲿ��L���
���3�߳0�k�������k٣����۶�g&���4*� 10,��������v�!O���[�^��Ǹ������5�O�@��ff��P�Z���D�s���s�瘦 Z
t뗊t�.E�18{C�׹����jA�p���Ja��]�f�#�}X�]�b�N=�D�쮣�'�Z�E�K�{�7��{�����-�
_�AX�72y`���]�%4cv�AX��Y�{#��ퟷf9Fo���7D�K\8��Cæ��C�E����DXjۏ�Sو���׆+�`����U�*GR�@�F����Z{3;��]�f�"́��CL�ذ��"C.�M���q��J�YG��6\Q��	e�ڲ-]k�$[��7H�e �-B��$ŜC-��3!������.:L�n	�_�2��d]z�<��2A�3D��u��C��Q둹L�� 2�$&�TIF��ٌ�����^{T#���E�~v����F}�m`?���Ǫ̂�����'z*��ER|�4΍V�����E�*�jPki���A�������?�B�Ԫ����o�*�b�-�i`��rU2+$�?J�8Z>�!*0_Ŝ6�5�3gOr�S߅8��Qh�W��E�L��U)�+�Ʉh;��뮰�yXLR��u����7q߂	�
6��������@��M�8�[��Jm;V��!�mk�)&�&(���vq�q!�JҚh�#���]�Jex���^'����'t�@Z96����9&[3��'Μ�k>�ͦ=����⇾C�s=��p
n�9i����*�~��x!']�'؇�.
��F�T��v1��B0�s*�N1�:�ʖ��(W$D޾����ٻ�U:_��_��ǆ�^��x���D��LC�i3:��w2y3se
cH�C+Wi�����׹���0�����gN"S�}�jO���9)������h�Cl���&���t�e�3>	�'��-(��<�>��jN1f��+|}�>��&��s�b�
^��G�{�_��,�\�çQ�	�IZN������o���|q���O�V��t6�� /Ό�[e��#7Ec`��&\��*�-�j��v�V9dh=������ա#C�ʃJm�$5W6��]�ad�	�J��F����6q�=�&1��������m��/���~b�y�:�Td
��Qdl�p�M��H(��1vZT�NI.q�� #C*�nıD����d��� ��d9�Ў�/ːH�O��J?2;���J@�z�4pJʁajQ�K3Sl,�Df���e�/V�r��y]����r�'*e��?s��-	�r/�#z�#xL�If(F%>͌�=څ�+�T�6`�<	���b���N�*g�S��-�T���pŸ�/[�ܵ����X���O_�![(*]kG�:y��Gx�6<ȓB�����C���f�C�$������ ?����:0#�n�sYԝe�#$T�7��m��W�2ju@Ѡ$ෝ�����$O��o�ӛ�&@�c�G̚vW9��7T�okәu<�l��q�i'Ieo(���+7�_`-*F���/�~Ǒa}���C�g ӓi�>B�T�?u��i��3ؔ60����a�w�{ť�B�m	g%�������n9����v(0���Tz��\Y3C���O�\�-�Z���b�i��@�����v*�L
G��������X�6
s^�����ׄ2ג�e7F!&��ɯ{��p��g^��U�;�-+�#X�7�R�N���ҿhl�u����K�����9ǝ*���z���/��_B�O`{�X�|}tc�ׂ���k���m���zF�)�H�C�L��-��7g�Y�����Ӯ�x��}v��hgI4��$��'(\q��/�"���1d�k���<�f���F 3ԍ����>l��v"���FO�gj����^*e��=c�6uX����@'�AՃ�EN��v9���-��S��<,2��'tׅ����.Q
��A��"؂��(��or��cbb�Jz��������Qa�
eU/�~�.�=���C_8a�?��עN83�~S����vҤ �^��uJ^Q�ăvMg\k�)�ٿ�CKƾC��4�V$�xi�*�`A(�1���G	s6�~�LϞQ�-q����庋��$l	^q��j\����ܵ��b[�� KײSe+�Tbjc���V8�z�r�5#l޺�D�ˡ�0Y�s�2�\=��9&�DWwt?t͗�z��\���Si��q<��Lu�Vw��UZ�������x�����x`ć-�L�9�O���'���!0��{sV�/��kO)"h
�?&JĜ����(v����q�\��~��k��95!͹5Z�k��eg��;��%�&v���Z��Q��fM%Q�Ue�O�v&������`��M�9p�t��O�t���Z���$�0Qە���a��O9�{߯D{^6 H6�����L��}XM�Jf�9 (x�,�3�b
�������ڟ�}H����*�Z������^�o;w-�O�n���D�~�0���\NR7%�>cC <�?�ߤ�׵9�q�ӄ�+dZ�9}�1�T6��7bG!_��ItQ�ť�Sn���C�zj5�0}��;�*�T\C��#��9�j'�3�6�?@�bhd^�I��A�/�*ӎ����t�6]\ͮ"���޻�gLj�/-�O-_MN�����PO��:�E�@�Uy+U�=E���?1p���L@�0�g�-��!�Yg�R0� 4B ���M8�����c#�n�bn0��O�ǿ3rn7�ì��Q8��`����C6z}���r���D��r28���d���Ot�2�8�I�r�27i*-�/Fkn{j&6�%�M/��Mf�pB�I	$9�ƣ[��*�N-�ɷ��d��V��VN�@�)]�/���ϱ��b�?�zع�J�=s �6�K9��rpv�BX'j�Q-�N�Q ��k
������
���9.�=�6IAyep�_�Z�
�zЖ_ՉixI �/�7&�O8�׏��?Jr�k�W�T��R�>��@�|.����@R�c��"-&�]0�{ҖP�E�p�	�o���$S+�=ٱ�PI��͊��M��r���;���8���O1~�/ay!L]��ʤ�f��@� �*g3�}V
�:�G�AX#҂�Tüy��]d�i�s�.��>W����u�a�ݕb�$@���ڿ)p/*�Պb�J�_TlNxd�8�B�5s+�b�q1�d
ޝ�A� �NO���J��FC"2G'���~���"2Vv������3gޣ�H�����~yq U�*K-d�32������������+ �w�ͦ~���e���X�6��z/k��T7�T�$��ӗC�0c���U�Kw�Uc�+ӧT_o!��'�$��Ƿs�ee�0<��uX��.�o���r1k"{���d�`���b̸�rv�K�l+U�{75�S��ޙP�\(O��#�7Ѐ�G8~(H':��\.�7��[(R�;��k�
��;���z��ŕ:6�bE6�6U�"k��M0��N����u?���e��_&M4�ꋢ��hd�.|6��J
�$���g�n͉��@7�~��8�3�|[&�zk�1���߰ςҴ?���~����q����
aP���:�6���v�6ww\�Cj�Uވ�Y���!�L�oeF~[W�$��5��;n�RS�<$�m���+\��O�k,��[�ǰ�M�0Aߔ��=J��J��1�ٕ4�c)w ���v�:hW��N����D�u8'P\~Z��}�=�Z9;3t���!=�Ka�} ���D\<�+G�H��b�r��mYCo�;N�n��[��L㋹�Y�{���n���%"��\
�NL[o����r7S�3�l��k���F�آ<�AV/�2~�}:��6�?�3���ъ�˝�D�HZ���=�<�E=�(Is_E�oP�П਒�;C����'l����d�"��SI��
�ݫ�*�H$�7Za�sCtN���8^B1����!�~��M_${�:��o�.���k�bU����D��0�	&o%!��ݰ ��-|c�1�h���M8_���"5m�*���#�!�� p�*� B»�ħj��f�t���H���j�1�X~m�e�s����ʾ1J::?�F�����O��|�Q��5���{$��;h4��y��'�=hW�����פY[�U�S)��Y�A�"w��u������ۧ�Ӱ��iP��I�5o�|Y��P�dsdtՎ�Mϊq�=t�����D!�ƨ/����W�GK�w�mx�P/%�{A��f��eB$Ȝ�D5����y�zȤ��������'��r.ǁ��R�������V���-r��#[Oes����|�e$4��/}($��k2?������G���CV��#uD/#��t��4Qo��"�4�g�5�1\�z��?�՟�C\�sUY����1��"�ü��;����Ƕ隋�38��F�K㲦�a�:n���)٨�^�%��5�ɥ��Wj����X�wȻ��j��5��� ٻ�=�/3n1oe#����ǐ#��{M�n�ʜ�,�s��$�f���&M�P��{������l֯}���5k�"�J���j��ן���l9�p����umW�T�n���eIy	-�z|ᣯe~?W� �x���j�$>�3d����C��#��Ǔ�D;���N���\�M8$�K,�i�i[g@3U�������OՀ�H&yy�8��}��er�G+��9#�����������'����x`ν�NK�CB�ڝ���I���/�rIy g�"?݀����E*)�u/������&���WE���(�JV�/m�HĴk�{|��WgW���S��p���@J�yѺ���t�����qz��祑�n�4P��0p1�;W�[��џ���QO[��!Ɋ%&�ƥ�El6A;�̀��b$��L"���˄�Q�4+��A�� �X�d�V=W���Z���h�q��"���2oe|`8��H�LgK.V���f �q����M#���E�ϭ�xmYƱ��^�H�M�H��o]4�����ǯ�+��:@/
��G�,�S�h��w%gז���r︋�tz+U��K֐>��l��'XW��#)8Ԛ�\�ş~_Z!����NϽ��q�*����voi�6�m�g���ǴKœ������c�^���M��J�wmk|kWAA����"�$��l-��;=o�pC
�^�����0L���E�)�9�[;뗐�0F�F�I:\��)xiW�ҽ�N����ոQ�A��d�y��.��ŉ���HkS���1-�Js�D���?i ���
O�:�����j/�ɝs�;�-ߝ�V���hb?������G�����)���^m�A2j��K4���dbf���M�!�\��ڌ����PC�?-����g�#=��C���'rxW�oma�	����n ,!a�����l4���73�PB&)����1�S���m�&D��i5i�dx�/���f��������ċ�r'K^�5�������]�E�j��8�̓�ڐ�*��ذYx?'��=Z4�'ݿf`�*+��s������Q>�f)U疄�S����)��՞���H�!Sk��Ŵ��$�i����E9�a��	�R��������i�]���gvE����9[;� �Gd��q���e�������|��#Y�]�&b�����$R�I���n�)����k(Ѭ�ƛd��d-�)�P����"g4�=oS��'�H�raF�e���\���')�Dm�Al?�8�>���&�7řɽ�X�Z��xm�\20�핿�w_1�o�s6|YZ�u&��򹺔s�9*�6_���K�/�q����N �g6��2���v[�$Y��S��FIn��9OF�>��4a��0�B����j}����L��&��h�R-�afO�{�ɦ�e�m���vˠ�I�L���[��_6s yO����`���H�p%�s��ۥ��T�I7;���?��4����St��ڿ��/��S�`�ߖ�.�?�' ?��|\	��N$�,� �Fі8�N����k3�\Rn(N����f��qS�����f������Vi(�rnh7�˖3n�&�������{�1�gǧ��5R��գ矟kN�͜J��m��|�d��,�)�<�SZ��f{~X��6	s��Z$�gKҍ���?R�z��@��ޖKu�K(����*����ϫY�E_:I}���n���@�~�T�8�5��̀���� ̨}��C]��Ƿ�>n��T����Gd�Q�Q����Ȁ���_�#ix�n���-�g���܈�:�_�=!H��C�D��{?�8�����{�=��{0���D3�� �0)�F3��jx������%�/���qA��sJ�"ը4E�z?'��o���h�bn;�܅���J@��r��j�H/��b�^�v�z"��(�ۄMu?;�M�xۛr�8�D�,"��{��.���r��u��:����Y,ZtB�O��M�:�R!���SB�^1��������YcOQ���0?�<<�>��0��OL����vQbX�A���q��o�}�?C���n��<�Ф�
�_�s���D@sgO��4����lM���H>3#�������"�\�Qu�iG/{X�Rf��:�E!g�b�%� W�����Gc.��NQ��j*��&��zj�U�Ӵ��KT����!�������}�0�ǉ��V���7���{��O:4x�#%�ӎ��~H0��W>~��PrX���SXU�JY5�:m�D�WP]8��YM� ����?�3�����7�U�ˇR���7�	��|�b�K����0��Ć��x��?_Zk�e��B����辄�� :�aD���Q��4i�<�0CVX|L�_i�����0�0�F����R.�y��5�ϥ�%�-��o�,m�O��@�k�k���8̝.�Q9.�\�k`u�mj�R��H�b�1�;��9ٟ��[yv�_E]��`p����i��` �)׆Sc�s:��󍵯���KT��L�00p��\��(И�˕].ߵ��?w*��gP�@�,-�@`��+�Ι��.��Yx+�V�fk���fN�賶�f>#
��o��g�"��ŏ�0��v��z���C�J�K�4b�+�UUJ����]��-��)6�7��S΅v��zۚ��{�?;���zW���>��^��(?��+�Dǩ�U�&Č�C����nx=KE=�^�
S��}i�iy���n���+\4�:t�HA��Cߠ(+#��r�?%���$ߟ�����HvO�۶	%.q��+��� X ��U@}���x\§EՍ������=��6M�q���:Om�&�XVJ��7����cߝ�����`���u�t�J�mǫ��ɶ	��O�8�j6��5539�u_vd���W�nͿv�<����K�g>e-m8z�l��ۉ-}Go��[[��lm��e�2�	�Ot��@���K�	̺����A�h~��85Af",T.0�0�:0è�'�pG��������(ZL,�`a��e�IAK��3��3�qaB���wb���
��$�����:��& PK   oI�Xډ�'��   �  /   images/9b01e4e0-397a-41ff-a8da-0d69e8cd9d76.jpg�gTS_�>��ş%@hQ�t(D@B'"RB� �(R�@���zM$TARCB���gf�����0k�z��y��{�s�}�}]���9���x 8��u����1�cǏ;�}����In��<��	�]�(�' p�
��%�����熨H$tU����-�8H�_A؎?�}��7��K���?�p�gg�u �y6��lG��+ 6 ��;�߁r�8��[��������ǿ^���n��\׎�޾w�����no�����߸�y���y#���VR�V=����������z���: 8���wx�� V�����?����=4��K�I�gk�-�$rPw�ꯓ�?D�X��ۮNL��}��?|f��z���C[��_��?/AϊX��ھfy6�*��عKM���6>�p�G}ޭwI�
e�v��{ѓ������vdK-S$4��ɪ~�ӧ^�g�e`��?-GՓr��.1#&�KO���� �&¡;�;χ,D��;��їwhk��)�g���:$�;�/�V^*xa�g�Q�Ta�5#j��M�/'^ؑ�t��"�����4�K^%���ꂽn�/�/�T��	�R
�.��%��[����$���D	na�"p���.�`��R��w	^tU�ڿbЃ��q�p�胾��s�_�UvƝ�]��tмu��[����m�k	�@�����v���]2�N6�ݧ�L�B��#���i�Z�����#�{5�fs0�@ӽqL�y]�lη&�����'�=�p�����#��� *?K�r�e����{������侍����#����ʭ��T����滗���&����޿��l)[ye�a���c���wN1���f�<�0��p��x	��Y�~g��x�K`�X���� '^z�[�O���Ѧ�ȽY�;Cbjmg��^z���ߧF)�6�u����u�����4,_I?!j�o�<�8e�mS�w��r5�y+ �i�;��Ƹ�!/��u��] �W<�|�k_C(�ӿ����i>��y�rT�j�Z�Y9|4̛�Id�2��?�n��aE��a�s������j;�n����@�_퓚��!�Ր0�8�!�t�0���z�5���3qlm�����!����l��-q�5�ӋA�MX�T�H�K���� /Uo�?ը�N	T��!"(xe���Bfta3�!�<9����u%�h�r���&�'��GY(���^�d��[G�և��k.��`��}�D��I��r_�����^�_dC9	G�Hl
���r,��T���'�ZE�c�~}2v~��AW{ГI&�1��ћ;in��7DW�P.�)���B	�b��_	���|�������문��|�r���� 29�-i]J
��"�A�d^}j��^�9 ��n�� ~�I�G��]��w�u�ZH�V�ƮF��?�f�{���\��xݒ�E�?�P���Οb0b<��.~J�,��q:�ؑ��^IW�^ۓ�񬅙N6?�&B�=�@�߽k��l/g�LłMT�����ꏫr���}{(��v@�M�/b�-�?��k�#u^�Y���Y����G��}�x0��y����WF��o\7�Qoݐ����ȷ!�K�ߊ<{�;c$%��+����t�_��P�<�&��C����1���U (�:���L}��,��7�YR�P����I|�{��k� ғ�P-w�wg�4�2Q)���dŃSr{�&��J����?R�6m�K(Ii|�2�7 6�7�.�U^�2�q1g�e�z)������C(� d��	��H�G����F&{��4o�d���s��Q����t���Ue2�=��!�(%����ٺ/Z؁ �R��=�.o��'`�|�yT�KJ_V�JFYg?�����}�<u�Au�X1���_�(:5rJ�/�M���pN���z]�l`ש+�?�w/X-z1�>5�,��0'�d�hf3+��P��ؔم�?
ا)�vANV}c���(�W�2X���-�,o-�'�l������&!V��P��O���V�fi<��D�i�H�/��sf��E�D�j�̣��hY#<g�&x��>電��+	���d�&^����>:<�q�@���_L���q9�AӜ-�R	�Ύ`Q�;G��j�Ҷ��2���R�ItĲi�c㝼�I��8�����,�>�c@u��b�+(��?����,pݫ����Z��+��	r9�,7��1ζ�.���:��7�̎;���B���/w�PDq}(��+__H�=�3pq��ms������B�Q�X��Nf;���_K�繝���x���#��]���������׵ի�<eVAE?kˌ4=�Y�J�)7��u�R�<0#6��+�ۣE��иV��MY5����M8q\�ti�Ъ�*��Q�߹鎗:�J�7�����8��Y�V����q �>s3	0�ދ��#V��;S��?�@r^��?\O��@Nd����9�=+���t��\�84���}��Ϯ�f�J�k�#@S�GLqh���6����}QA|Pa_"c%��T�xi.�R� 51[��/�F ȧy�ob:��ϸ��
�Oҥ���\�(�K�	1���*ʹ{OI?	ⳛibՎ��)�G8�E$Y��i4@��+�	�V	�(g��F.Lr��\k�� P�k�IX�*ӛ>�n��D��G��'K֡UE��gޤ�d�D�Ӌ���m��ʈ�|������v�m�m
::���h��0��jθ��[-W�R$��;�i�}� CK*g1��X��iQ,N>��b��(ϊpT�Ħ�W6�Q�Q�oē'K�����$�t@��F�x+<�Nr�K�"��4��|�%���r����}:�����d���~�l�%�<0]�V���mb��b��%����w�/p����;>?�*�{͊�
����u��Ȃ����߹\��3�ɉ B��e�E���%�JZ���G!O��u�^�6��$\s��k2��e�ו��6�.$�.�d5�#�|��;u}:�=������>��ZeÃ9m�Mv�������yj����k;�Az؜_3�U����_���4��$~W`�f�n�e�dxw�x6��a�N'T�~�3�¬�a̷Z��D�r��Az�U�ZA����V�m���3�Y�4m�a|B�.����:��:����P����U��v�Q_ZJ�J�(:VZ�v\X2r@���9���i	��O��K��p̥�l�kV7�|~��_ˍM�_ָ�2�J�D���?�������G��i9>_������)���R�y��r{��cn9۴�\��A����K2��PH|tҟ�5��L�����������[ps�|l�8|�jQ�w�[���W	,�X\��������tk�����h��}R���t[y�`�m\���9�~ ����\ʜ~x�35���ѩ,T�/���-�pG5��	�x�a�ph@��S��TE3ʂ��u*[�ë�T)��;�T�&c�T>��%n	Bv��O,�V����G۳��]{F[�?�����N��R4�]ɬ�!�g�ƈfɸ��`���`ш�����t���.4�P�=5��zB��ߩ:��s�ɢ��R>ц-I��Q.\gE�QmqZ�E����k��)�-��|��k�Vˡ�5س�b���W�C���.w�������]�=6I�ؚ�t�n�J����l�1Q�87~`�� Q��1�<�S�̷�<�IA8� �^p����U��(<H^��h0��+	+���6F�ʀ��#r�$֔���n;���dfx����{9��!٧|��>�t�;b�G�����ߧ�ߊ�ܼ�[��&tmB�i�@�,��H�!m]�]eW=w�`�h���&���F������Na��ON9�&x�:��0�64�mzsxZ}U�c���q�޽LX����)��{sx<�Q���f(������&4
��)�&�{����`�5����)�q�ӎ�7���&�L+C��X�n8�^�^���M�,)���$�O��H�S�����<���~�W`v���k�*M�D4�D�ކ��_�W��	(��i��\��V���
��қز�~��]��R�Z�
�1����<�Rk��$ఁ�O�n�!������/ I;�|��p��)�-˺S�i���'Tp\���R��7�L�:�޻�+F��y��A��<�+��ʨT��y�	����U��p+�-�C���N_��m-�#-�Ӌ�L�q�2!�"v3�,g5�V:}�ӄ�� x~�e�<wL�(�E��%p�Ҽ�9*ѽ`;#��р�Z^����3��6�����on��:jw�o�G$�h�A-X&��40�C�
F��]J�+��~o�T���w��FBn����/�����̥K�h"3|�~ ��)�1���d�2�����E϶o'��R����=�H������G�ׂp0G���ut��r�:���^'E�-�6AXgaf����(�����-�A���ۊh��R?z��#|e��v<��4�6p�3)�؈SW��\�A��`�.{�"I�n�AR���/���w�蛻 r��U�Ee�OqY�����S)���8Y3c�y[M!��@];�p��`f������BύH 6�E�[��Ӷ���H�y���o���E�K�Y>_�M����XY�~rA�����8?������6*�F�/0��{ؘ�����g�F:asX!+r�P���c�֌'��wds�S-��)9�t֜�!X?�Y"I�Y!u!Ѐ��L�f�+7T���Y�g���ˮ�9���l�	S��ߡ��ʞ�z�4�hX=����DL��ۏ�n�՚�B��H����Py��H�j�+�0����M�����0�ōGɏ��1��=��#%{*���*�x�w��X"�|I�)i���I��晼����#@��XH�*g��^e�*�I�ں��qzaj����_W9�k�;��I����WnV���m���d�y7��HS�R^OJ�v��˕y�U��-�B[��לƾ�*/�/�Ӵܓ5�#n�r������(�;���u6�!Q��I����e���.�,��N�r����d�ޖM��X�� e��d�џ\!�PK�� �Fr0M����!�u XA��h9����F������.QS�370箛;�/�x�%���;եC�,�&j>�n�E�N4F�n�c=Z��z<>m�7���u�m;wl�	����N�������<���n�3Ns�Y�S���@Ujd����-^�ӂ*#�����c�g�2��Eq\��t|��*�FKzĬL���/W��tO��ί����n���`�J�~a��E���_�20x,�٪��5�O��֘-�<"�������~��ҽ�S��c��@���z�]]�wj�d�Tn�P���&�;m|�[���������K/:Fu���>-*�t+���V\%�����ַ@4�E�=Ys�1��B�=Bs%)*�)��P�󐲉T��-C�͔e%���������].� �G#�����Ӯ�d�PX�L���/ا<��?�WW�X���˒��b�j�A��j�[��i��r�H=��W�{�SN����$�,ƨ�~�kӏ��uo6Կil��|,Κ�aDQ��J��Y6�%�FMh�iFQn���of�=�q���Դ�*P(��uEt������@װ9������)m�č�kK�7�2 ��߅t�&Zb��qg~ɯ����.'F�!�U���6�я�8V�5�RQ/vf������zb��6ӵ�5G��'8%��Xʿ�:tK6���-,,Ձ�w��W7S��H���=�6j=,��w�Ӳ�S��T_4�N�w�
������ؒǜ�{˜��f�;�� A�i����*��7�)>��$=і�E�/݊5Q'����G�0��7�kw�7�e}ڞ��d�
�-�j��re�ne����Q��k�{�q���N�t���1�p滨�	z�0���q$��uQQ8�l8�_߄�/�VXR�u0l����>�Q8�'��ﱫ1�~����k)�}��
M�i\��*k��2����!I9���]da��� h.�l�Z1\$��U��>�UE���f���ᆜ#��y�O"�Щ)�`�AL�����߳�6���T>�j��>�F����lE�Ms%&�r�S�7�1�^%����1C�_Ƶ)?��w2�e��=�s��=*�A����QB�8�g��D��s��LL��N&o�����ɊMI,�~m��W�s���[P��Z�K(QL�ȷ/C�C�#Ǿ\c�HL��g�G�Blz�&y`j���Qu`�����9(Ñ@�����Ъ8ù�l[�[;���L9sg����@����GA�a�=��l�C}BG���7�a���Z���a�Ӕ�,���l��`�|CB�a��aG��^z`���O���=ن���#_\,9���f��'#����jx�M��/�Mi�7u?��q/�[η?O��Ѣ����L˜QU����w[o��h K�K�4��'��-t;M�8KL-F5jl���EF_$�R��?��o�H�Ǎ�C�8��!R����C��s\��hJ��H���_g�IJ�Gw�f\�no"Wc�BL�5~�oF䅑��~
�#&ד�D@�ݑ¯��6Fm
�^jy�&m�2a=w�,�1n5M�㑑��*Y
����YA�u<Q�mC�<o��0z:*�(��|7��`kv��k���N�� a��4���7�;�DD8��f���>�a���rc���J��# V���̵R�85`w�H����Wt�Ө}=�	������)D��l��O��c�#�7�gg�N��&��w�EzD3At�V�r��4^~;��p%~����=���@x,#:��.�V�*�s�-�nH����B[}v�5�.��\�U��[]���p2ݬ�~�����ڕA��i"9�q{����u%+�������O6~�A45~�"z��w��9е������{��!��鬫�������v�E��M���a���B_n����<t��"�O:$�s�h��{i.�<�X�s�ω�[|��NmȢ}�,OX�� ˶.Ix��j�(R�π_P�f,Ӏ�]�ӎ�{>�.|s�Br�8�e�_�tIr�:v'��r'\o��`������:�M��I0�@ �?���G��m�,��do��=Zr��Oy_�ו����Zc"V��",��ƨ�+�z�:JX���O�u����G�7@�$�tB����1��[a^�e�)�w��(�� � y��6zE��1�|�W��"�����ɧ�nUC4��:��u�<df��<�[f]��"��t\��v���7�9�\��$I@� ��saA���I�zً�����K	�O�f��&�tL��.�E��}�vz��Sx����JI��(�wU���4���_������p�:	۷]���1~F�dJ�ޔ�?�&�S�W
�����;�lb�*�"�n؎_q�I�-�ik��^Y<�Q�:gM�\�E�,�W8�2)��;�*���"p��Ir����������lc�8%���!�«b�Sg�!ꦋ���L����t�r���ވ��q[%�ţ�(_��ም~�5��^.ӛ&���y~�<!Y񫴝�[b��{4���7�N��[o+���%aA�������TQ��g�aŷ�O�M��p��cx�����\�C|9Kx��ɕE����(�s�F	��6�A0F״��#RV��l���M۵��w��l�F�x�tT�c�j+�?�Ui�$'��!�/��d=�����C�4]���D8�~0	�>�Q��RW^�~����3U�7��Vrkh{KQ�bJ��ʢ7��S���a��$q����?��2�p�L��D�cя�
/a1�㟠&-�X��"���o��8N�)��Ͽ��q�< t����46~��,R��"�4�_�B�@�)4�	Co��j{K�C�۪F��� Q#�7����w���$/��efq�x��W�X)�@ߩ<���&E-�-lPS��9�!�n��t�Zd�L��اe�?)��P@�m/>��MkL��PZe:��e.��'��ѕ�U5O=��@>��!R�{8���$�W�!�l��}ɋ���]"�,��Ѡ��K�@�I�7nw�s�D�:�UOEbU�#�]g�����%���G������djL�c:Q���[�+S����Ǝس���Ϻd�Պѕ�Bs7nR����@Z��������9]��������d����F:���^����%nٞ������v��7t6HR�����A'B��Pt�+�{��7w'��Ú*��َ�	�vt�t�����~>k}Ww���%׹��,��Ȑ�E.�ԝ�LV|�ّ��+�Lw��:�������ݝ���(I�Dam����C!�k�2<	g���!i*� &�F}~A	�6�$�BT��>	;'���n澇�7��UG)�ӱ7���N����	��ή����0���o�%.0R-�qB�ʹ�uq�W�-�>N���P�-Lj���͎��2o4�04>��4b� ��m'\Mf�#��<#ܼ?r�&�:��]���3�a蜑�Z�u����Ɋ��;�H���_��*^��"��W�����8�-�m߈�lO�)O�,��'C����-'RIJ��d�s�M+<�L��7C���c�"�u
�LFdj�w��=�ßɀ����.�n<�����^�`�����^=Jb�Gy���M�O����$^��J�Ҕ�~�E/�Y?:� ���d�To��0�6��+�k��_�dd�G��֢/��̑o�ݢz����~��i���M ����{�RH*�K-�ޭ3�mUP�6�z�x�<���J\hvK�ђd<�~��,H���C_�5M޻�s@��f����Y[+�~�d)]�AgJ�Ms���%��f����m��;G#@{��*F�l[ͤD9]�ӛ((�Ƕes�B����ee�g�JN��wP/{ժ��߉��y���������H_��y�	��J#jc��Ϟ-5�u���N�G�)�i;6�?Y޹Y���r&t��#����B���Rn��(B��hu�\���40���g�HVt���g����%PZ��(H�r�@���M>H�r�z��}U�rP�8���G�!���b��j�;�#@Cye!v��Yl;�v�� ����=?�u��mҭ�kk��U'KuD����>�i<�����C��"�:c(��)EM���eߋZy���c5m*CQ��l($>HgW������8�]P��p��"�zT�I��)�^ ��|x6uh$����䞾91��"��)�B����A��ZYqDP��sK����2z���	��,���<ݪ3���>d�^�V��e������7 ;�Y��uܐ��?U��gtfÅ튏f^�C�R��2ˣ��&�]�+�j�*_̝Q�ڞ.*��٨qTJk�3�r�e�ʊQߗ�\�M�?�Z%)f�� �@�Xr��X���b!E4��Ӊn��r��\����Uz��M۔�aS�K*jN��n�Tԝٯ���E��!�p��W焯̅��=	��2~
����2�� Z��]����7�E�흷�Q:9S�>Ҵ��?շ��(U��]uh	�6wq���Wz33�S��2xt�2Co:oGᡕ��y��sa��"�!�T[�7~����(�(���96�}5�{D*x+������������vm��ЃHm~&X>D޾!��f@:C.`�U({ � ��>CZǎ�%M��۳H��.Μ�r=�A���CjL�%��� y���v��x�`wx�����2�&�)b��NRגY\����xw���;Ȋb���p�6� ����ڙw[S����ἲx��D�y���ܕ��*/�mG�*��7��j���%K�$�;|��M�/�М��͗�&����S�����=����	q����ޕ4ϧ�o=>�g��S���@z�j�T3�M�j Xbb��ژN���e�u��$��}r��e�R8�+�S��~]�6� j��.����'�P:!@%�|�K���B'r*�R�f���> ##&��1׎=� Vx�D��7�@�z�A��W��KU�4�ǜ�N��[`?�%��f6t��9u�� z9bU�c���C��K��~"��^�!!�M�e}�IX���B"��k��l��3L�PP�[�%=���:^YѳOw��Y�����Z_�rU4���]rP�2�2�TG)�^�ߣ�\v[S�jߠ&��X�o�gT���%�����e��)��=�`j�^�U�3���I��. ��i�F��?� F4���QA*�%Y��-T��A�$�.>/M��'�0v�V��o�5y��et�i7���a�����tp3���U��e�yMpD9��6,��z{:kc������ܸ�Q���z�L���}��K>�e�ȎI}<K��}h�1B�m�*��۠�È�j�w��^z\r�*��]CJ�y��wa+����B�XH7;'��o5�O�6q��)��2���c\��]�\�c�S��x�nosxE���B�������f�G��R��*r;T�B4�Μt��+��U*?_ޖZW!~�����)U�pY���������S�����۱EM�n�1�m�O:`_��w�l�+�ϗ��!�;:�_i�K�٪�8�I�<[��1y���0
s���:NO9nc�I$0�e�Y�h��^S� �m�Xd�H3��$��,��37��9'�4T� �$��Wp�*���f*���<kc��h���1T I���j�S����<ހ�������C+��U/x
��;U�|6�
��/Z}��6�5��q�y�m2?EϪd��q^Xͧ/C���~�/��ǕQv��>2��au-��e�m�a2/$R]��5�t��VS7�_���L=/e�[�ژ�ѡA�}+�p�^�СP���+��gu���)��������VR���oͲ�����m�?5|���&�T�g���*�6Z��2�niN������eɚ�m<�>�`6��V����ۼ�*��ub�R����c�Ăڹ%�#�'����}��x{���39�iӘ���B�yko���&�|W)%��F�/�'=1�ww�Fcަפ��d �ڳ��Q���^�v�ts�Vϳ���$isE��S9Y�~�ϓ�2����7�PXzT��w}R0���.E\*���=�W��NV}���.(RVտ��ƓEk�q;�Oq���wʖ�����~�^W]���..庺��7��>@����UdrN�Nx��w�1k��0���=w�Wz.�������ס0���r������3clF	h������B�B�dq,
v �~ -#Ji�t��<�
m�/���-���zey,�m>ѓڶM����Rx�����x�X�r���f�������)NZH��?���r�hz��)=S�48d��1Z�2� Au���[�77����a�*�ʱ�"B{��pA&�=��q3X3ɬ:]U�9��IW����:��6��M"0sk�IpKO������ٺ�ir�?
sb��J÷'1/�J:�13�혭98��̱���U�]�I6�@����'Cɟ-o�t��c͚ĕ���K��	�[R+Os.x��#��T��wb�������b��>[&'�Y�/iCG���K�bG ����/�
*�"p����K�W�h�Z�%��S�����|��,��!���!!�t#����>�:2A�G�K��GP��	�(:�b�0�ѹGB�RH_�Ώ?W:���pR!�\u�%�[�"Ξ�[�U������S��]��Gx�h��3)��rs�+#c��D3�5���/ei`��5@�0(_����O�zK��j����m�G77=��l�P���/�g	�Uu��s����������סa��C�)m�x�5Q�Hxǆ�J���{N�qf�Nξ�z�,�#g�(���aR£�\����] F��d�2�-����2�N*!��he��`���a\����;*�	��Ш���vI��󚹏&�;���j2�~�|	�l��FW�(�w����[�u��F��|/�B�0$�dP�8��W:����n\{^�up"�������?�EG�N�����=���3��x�p���U���ƕ�;u�����{h�]��\8q��U�c�U�j�e�=m9c�,T?���=�|�}᥯k��/�E��{�x��V����# ��yb�n��H����q�_�6;H��ԙHwv����rFif�ȡ!��xE��ߢ�p�uXߣ��F}�b����b��Ċ��u��Q��e�lEɰ��֨	<3��`�u5�x����9������hBP�[H�ro�/s�
w��"��y��?;|���-��`��J(�(�+�yno�W��J*���P�b�w�����Ȉ��H�3a<<����kF7��5��±}a��<�� ������O�J��"6�)f�!����aU/�6����^��+@�	+$Y���*>׏�v��;�b��now���*cE��F�.�B�<����n#�j{$�ea�CH�֙V�i�j=�� n�q2'�b@M��w]u����<��og�>�	-:B����\��2l�!,���
2�F�S8$�u��:���N�P+O��B��nG��V��?�����!��I��;f��V��AH���+��:�J*�~���Vm��/@�DL�jxf�0F�,;�Bv�Jg�׍�;=�������Y�������i����'�����)�齞,�#@\
ֆ���uIT�8~���F�ml�/� t��%������dH'�M�L0��u3�i�g�S�@$��f�}$���Ȁ�nәX�%i-*��t9!|�_
�q�� '��[s�x�����~+���=62����$���W��������5or��E�X���	h����YbNd�#�|�u��g1!�遼y�\�BkZ��-�&5�+���2���ɚ\�Q������S����KXC1�!M�\w����3�i&�w�Q�^�&�����*FSy�=���tfʼn�%#cq�:�Z{C���@c	���G^�6�!�A�Nm��4�$��N�N��JEk�-RO����i��1����W ���-L��Ul�l��YN���"��!���d��R���b��3��Ҍ�ԡ�F�P�w���
z:�9B�wd2&f�e.����p�/=b������࣬���Iҳ�Z(Z�n���)&�ݮ�l��Glbc�/�@Ю�i�LE�� R���#�V����:��fEo�6��>���6�g_k����U�ĩ�,�8}��X<�:OO5x��qc�:Ik��4t����#JN�>���i��t�f��Iy�F�n�a~�����N�5��V4��7���Jxc�%�O�c@��e�7�b���k�ZE�hqL_��k�)m�+��\��\ҋ�� u�C��y��S(yNy���oB�"n�i�����JQ�'D��/���^(�[��Vj�6y2�5is#���|����(%�P!��.n7���}��o���c3���|lx���u��:bi�p��ek��$�2�(����m��$Gm-�����U�ܯ|�����ӻ����2My���P�X�W^�?�&����.����%r������N&�+���2��C��j�m¾�<�}����ED���9�_8�v7I�Ǡ��ALR���o!�#@�ɼ�RK.�Z��Ju
�l.�Bw|nB?RJ5�oȸ�2���=�;J57gۼ��-��	�����&���	L���%��L}ֺ��n!�u�=�x�VP�/cO`%�W:�'�̚��B��ʈPy��w
��9+ =M��2@�;ek;�{	e�#*GH��S~�D]��ּ2%�5�����7�)�y�),A�ա-�o����>�("���P��9�$�(���#��)��4����hܨ�  �q�-�!�F��1��Y����Z�'�1�9y���V�\>���Yڎ\�+��;���l~���6M)��>?#�����x���)�>�,_u��Iʎ�%��¸ ����f�����W%-�~RJgi�)��UGDrm��&�Io5�M % =IL������o��PR)3�&��*�J�h�c��T�Ǐ>�詍f�~j�ϙ�����)�ދւ�x�'��b!EC~�[Qz�e`)�������O{��>���*��w��n݈���K-V����l?9?���� �+��m�.*%�E�1�P�k�E?�>�f�R疯ߓ�ݳ�,G4T�2�,Ut�,4���|2̭�6�[���R�,���t�nHs4��v�T{��,�{С�4�Q�|up�ߕ�J�4�kf��_pZ;�Ӈ��'	���K��⍴����y���S�T��|�2�+��Y�+ȇqP�<�R��(����eY��2�� �t��Ls���My�x(�,[�=���z��41<b�� q!P��BO"K����ݘ�a:�sYoe�����ɻf{�Ӯ	U�j_�#\��R_?n4~�dY�R��y�՗p�$��&a���KZ� g�Q��.٤��"��#P����*�ޠ�/�4J��iB�SŃZ�������F1�ٺm�5�+�l73���R>&ʩ>����x���_����WQd��}Gѵ�=������I�x��Ds���8��ǲ?M��ز]B`�m���u�2o}�1x�ɴ8a��ݍZ�VO�V�}vm��yLx��uɨ|�Sm������8��9[��~�u���gI�����z+���w�J���P�
�����x��Y��~�`I<�0��+KwU��g���y���ׂA��,���}z)�c;����І���g�����C�'�u�k�＜��ӿ��=�D�9���O��i�[D�z�)쿧1�VS��Qǲ����?Yfc���Vqw�SƖJ�w':��4��<���*����)f���jy�������,�C[�*��Z�H��&�񃯾��������r�Ț�j[�ʯ?,M��Iై#�9�s=��٘�d8X+.5'�d���l��ʾo��L>'Wrh����*X�BT�XЩ�Tx����lZF��T��TANM#e�L������:�� ������~���#)Q2��EtW��:��#���u�����j��m^��w�����a_��� E�n��>���D�k���� �����έ��gk���1��(��(	V�k�m9��"�P�Sl��*!�α���z��5���$���|Nݯ��.�jӤuj�=k������}��Xfb���\<.�t>�^�)q�0��/��>h>k�,UX�#Lm���ψ��+3��{��'��4��.ƥ�A�{��<�k����@�6��/F!l�w��ypv�N%�݌?p`AM2�ilH������!-��{�wz1�O�u��7�����+�5�E��K�q�L�F �;iK��Eg e˨����#���V�
�y�n�%�$��_�g&H$�F�vp�3�яbb�]�&��1^;�TxR��{{F�*z�>ns�)�d���L��Y�Xe���QhR�T��%Q���6A��s�H-w���8�/տB����Z�+M�wd�$�w��M�47瀢�Z�#��I*��i�版����ۏ�:��,KX,��ͪ��7�Ʋ����P$u��B�u�F��c:t��(�K�����o�Viwv�!yY��͑���KǏW�-���L��f�B^8��L�yl���`%����mHv�����~N�S�#�O�K�ԅ?���rj����&Z�R_y,�}��>�d)��x� ���P���a�b��V��"l�PY�+�I�?����5hqmD���P[��p�X�je��Uꡝ+Ƅ���{��8u�v���9��u�-Ԃw��J;��$G�ͤ7���Uo6���s� �ט�����6zq���Pϔ
"��*�6�r��x��r�P���z�Q�S�5˩n�
BkuD,K{������ȕL����ͥ����1�E�[i�C#�7� �f}��|��ڴ	�$پáC&����4���YWU^�5�?���i����f&GiP#%I�FV%����vE��!s��P����)���sD�v=��n_V~��F����ŹD���uG��"}���$HeSU;��2ۡ4ن�ih��e����Y`�*y���D���K+�
�'�����.����:3��4�~@���!�5�?���Of��^r"L�o���W���� �* �Ҥ+��r	�B�T@-RB�(UJ�!���J�$ �"���!��s�����~1o�5�����f���5l�V�?�)�F�q���i�z�%F��rr?�ThZ�Sh�^�)�]i;;M�^�v��0�2Ǔ33��6�υ�a���C"$jC!6�����S&��~��d��hd~������!�!it�ko.��X�h�Z�=��m�|x�g�l�?�&`,����߿N 	�{��Y:1A�}�����'��A��-�+�@�Q:B��L{��s/���	 ��[N��t��_�L���iV�M8'�:�:U�I��<2�x)�e�lw���	a34z���A8ỏ#�����F^�?��<��_ �2�ͭ��FXpPZ#Rˎ���A]��lg![Va��]�=D�:�6�xuu�4c�aD��vY�,�*JՔ��!k{���UZ�(Q�4��s�Z�=
eQ�0���l1���Rd��u#�tY�k�;�G&nY+�t�b���#�e�Q99�tiQ]�o���YsԼ(�g��j&Ч`��n氐��F&�y�n�5����G4�i�&#�� ��KW���B�����w;��[n��8�iѺvl�?�wä�?��k�z��	;x�ѻ���S�vQ�m�$�*�a{)���z���!�M���5f����뫩XrL���{���
����T,�l8��6z��"��3��LwS!-��fo<VO�q��z:�k�E�]mT�V���"����:|g�M|����#�������F�%S���
iw�\y0�נ�U/a�?�}:n�;։�{ĩX��{�]�8G��a8X�����p�:�f��k�v"q��&��I�02�݆�%������������#O.����=����,���P]��Z&JI�� Շi��M���q�T*d\z�c�V<z���7�Z΋�m���q]:ǯ�yo�%�QI��1R7�r8�|�i+�*�;C�2\x]���%��ֲ���U�к0�hQ�=vθ�p%rHu�=�}����,��C\�}|\��E����#:�Ÿ\
�1�1PȻ�8{d�~��E#)�u=$�:}z"�@�mZ����U��v�*���O���%��og��w����-g���i�z�=p$)EI�Q��L�4�T�M����������0.dF�� ��9r�|���1:�|�x�����/��D Z�V���_�XZ^���B�0®4Z�h�}�>BG��䁇C8��K�g��|�u� ��l�Q��,!;���,�[������鑬�gI�XMԖ
ԟ�}��{�RR{�X���0�~��6`!�0����?�kl.�^^P�"�c��J�d�O H����d�ܬ��/��ï��8�<������)����%�>�u^rj\��г����������������f��xT�?/�V�a"{)�^����{%E�N@�-Pr�T�PυU�B��7Q)��ge���x!�����/��G�o�ȸ�=V�x�F�䴝%����T���8*�.�H|�H���RX�92���0(�O�����{�A-� j�c��A�E�=����N�UǯI-{9}tQn����(��i�����L�q`�q4�?������pm�V����r֎�ʻ۬�H�!�̈́�*μ9bR��\7�%�
�x2Ic׶*��I=ؓ��8Q3�an��UK���!��.I<"x�C�Uʵ��b�����X'��l�{��6hp�?n��$GS+�M��SjɽZ��ŕWKuO��{�ԚV�����ʝ{�Ш 5�!�ў1ޡ=nt`c���ǻ��/��)!��E�AuSFz���>y]�ߊu��o���ő�呁P��(^~����KXdz��~�(�^9�J�C��%ʈ>���e�@��	�콗��4��\儫S��e���濷Crq�0�kQ��ѭ�}k������X�9�R�M�I��ʂ�Y��u���r��E�r&&X���}f�r���E� �Y�W�.n?l�����[�!�r�k�fk��L�A��$P��fę��)A��ֹ!�w@��>Cn�oz���ŊY�		�(����z��:j9�^���)1";�a�`��fe�3�;�H6�`|5�8�Y���q���H#���'W�Z�פg�(!��0P��-:���b#���@��2Z���ߩ�j����eTH26�;hu��y��0K�|;x��
���e�8i�{�ɶ/�6L����|0�����K焩��J�����䜍n��i�H=�Q��衧οH��Wn�_�t�J��v�ǋ�7GO$#� +�ft�ǯ)�[ʽ�f�k3�H���
)�ö!׉�M�>�-����]߷s�.U���ͮ���J&�HB��~������-�j�60$:G�X�{�$<��8\T�ޙ���`l)�i�yH�o�:�Vopi<��44�A��b�I�o["��#n�ϙ pd@������n�J|�)�`^߯��2'}K���2i���.��A��%+_39�ɜ��L�o��sN�9r'h�kf!~I����?v���1*&�~C�MJqB�ÿ�!��gn�����n��R�kvo8M�*��'r���0�<o=!�Y*�;�Fu���ǖ��m;tu����/ueZP�
����y�#�>��*��Sj�|��b�b�19��ᗽ7ʔ|{�4�V6���*B2�ʌzb`,o���_Y��>��RW<UAxd�&��/��8/غ������������¡�PM�a�:���	�����ʁ�U�)6L+l��LUq-��~ղ2sc�N��(��zw���a]R��ѩdO'?�w2��3	�)���Lt����,�4�lƗ��4d��C�����878գ��B�a�JS��-�I�jz��<U��s��hK�Ncν[5�72�I,Zh��baè��r�޼��_�I>��._9��6��ܰ���j9��<�z~�b��ܓ����%	:���X�[�h�5�iLk����,a�O88w1��ZY۪���|�k��o�yAT����tU`f��[5�.��aɰ����V~�;P)��uAZ��&��0F�_���؊=�����������r�I��b m�h��]9���#���˂ie�3c��Bߛ+Y5���r��;�j<r9�h:}wO/�j����Ve`Yo�q�60^u����U$n�7�T��|e�[��0ט���I+.2��.aq ��-$��>�?c��aS
n�T�������@T��X��:�ex��G\�q�Ey�@r�zdь�u���o9^u7|�c�RR�����j��OoJxO^�Z��p�4~ ���1=��l�d~2�B>������yc�Vv���s�?�����֤�Hs�cS��!�2*��}�"C�}���4m���M�)�g�ʢ��g;U��'�|h� D�>���^-��R�̒���]r*��U6?<�����`p��T-�d-:�$f��� s4�$>'[a��$�>���>��1ҪQ�^�q<�`
=�5C<���P !���ϐz`;2��+���a��.y3&B�'����}o�6g�@����M�c�1®(�d����$��E!�Hy�
�;����{���Q̺��������쬦(b��ڰL\�]ʷ��G��x�;:\&�h.
��YA���&� �5Mo�l��{`��k�>r�����E�z�W����Y0�}_���]�ܻ@�F{��W�cc��r�P)
�������吚pw Kz8�B�ĵ8$�UsH�����
��JB_��p�YyvQ#3γc�N�;��~T�YZ!~��,��3�P6���8�����;�I��Ҡ<�+����jO�>�s���{��/��!�����a7��l�*3x���B�R��*���OB������]Aߠ���k�7ˤ�H�
mt�>8d�m{Lx�e�se8Ǩ��*�2"L՗�ή-φQ@�]̿:eU4|�v7��o��Uw�U���^n	����f˦`��p�ڥ؇CTo�b'3�Ǝ��{C�r�Z�
v�@O��e��!�{�kf)ݞ�������'�:�A��ؤ�u:ϸŵd���ʰ�B�خ)cUt�C�NL��n��κgWX����5d���kMjL﨓�K�reMc�*1����R�H&�[�ʚm���^C�,1��?��X���J��gHX���7m��f#�b��c�|�1V���/���4%����c�1�r�O�B������n�`V��<�iR� �3$�Fǹ� �yJm�y����9��,��v�텗~��O����6g"t�~F��ܺ=�9p�����? 2U8�.M|o�<�Zz����>�͏�ew��3�,���e�_��u a��x��t	|�8��%*И�͒	Fի�?q����O��X. j����Qk��K��;���Ƶ*�y�o���޵�ߴ�Hn�C���G��)����ZXl@��	}`��i��Rz7��
��A�9	#��wދ����(x�M�|��֩�x܇68��%��[ 	C�/Vp�K�-�N��z�8Ȯ��L�~���L��k��O�	9?Λ�Un~�O|�]Uk����FY�#te��>�)sڴ"&;���\j��)��`������JSͱ���V`
K�\�R1��+2�x��������l����Z�����{Z��C��Hb��[���������t�������+	vq37��6?|�u�}��)�b����]���w��w�����C{���Ҧ�_�����޳k)ë-2�-d
]Kly�r����~�R�f����0�M�7z,@�q2�F���^�4M�L�RX��x!������z�8`����ϖ�5�@����;Q�F͈y�V؛�D����|�u�/�3����I��ˇ�o&��ۀ�y<�ӄ@;- ���
0�<�O���9���TS�jƯ��8�ei������4��hJ��ܙF9e/���?J��%�����b[R<7V�e1����ۧ�㥗Sb�8�Q�PW`�D�-s�Ԡ���=p�w���i4q<��،̰<R�PDd��r�)���dбЗt����O��q�K�"��ov�R�UA��'�l�#�C*��ź�� e�ɶ$�������	�˔:�ɚ4
���`*�'��75��e�+�����CbZ��Ҭ�����ݖ~��V0��*Cy���Od���΂�W��Lp���S���Xa-��3�)���fz<+.�^@�о)��ؖ�eF��9HŢ�%#�n�M���sJ��_�/�_�p
E {���>7%-��\�+�n=I�D�3�"��m��� ʒw�y5�r��/-����t@�}f���k^��g�H��_|��.��^gI�~�g���A�ɿ>$7�'N��=��������k٭L��ѡ61@�^�/h �hg���o�8��;��HW��x�(X�ùP\h����^ɐ��'>4$�����^v#��n`U�Vq����Ҿ���4�|"A-du� ����D��֮L<�]����P���)�W�Ȗ�V�Q���̈́��|M}�f�[l0�:��>�$�M�5):VAXb���kNm���.�C�s.U����@.�/��֥�&�-��M�)\U��f��i	��$Ex��I��_�_\*�R,;o���1�� n;�/Y��=?�g����s�
��w�Y5C�7��@q@8�c�Z��G����ފ�fq���؋�=F��Tzudj�۵��t{/���>��+����6+�,C���׌0��^�NM^��ƅC.D�up嶌�g��w|�a�@4:�)Gms����>�Hz�<F�1a�BU�_�0M����7�j�Ҝ��o�2HY�֡	<�M8�������I�. ՝�+�I�ih43��ԫ�?��(C|�Ֆ9̽�^��R X���|�6��� �6e����K���'ky�G����8Aw��;��^�� >|�^S	��H@����3�s(��b[|;k�IO;n�2S���}��O�5��zy�9���|��h��MȞ�Nsbk��y�sWF-����jx��g|� �#���
2f�P���fM F�ݴĉ��݇���M��ML���C����IU����E�<�z�x�fy?����8Ƿ�L0�8�v<R����\�q(�i����b�;����t��Zz����g�̝��A�q0��M�u�ZNy��0���o����S�\+$;7�ܳiJ��z8�����S厲��f�L^��|�k�I���f��|�W��\���R��SІq��� x#����'˨fc���ظ�a����_���4<Y�A�/�K����9��D`5�穥�8�ux��#�_��?��yH��Ӿ]�-ܸ}1�gb��� '�w3�Z��УAW�/X=Y\$��n��S�3rH��}T���@���1�܃{�J߇�`��.�Y/�����~᧓���<6%�/uD^A����c��D��xʼ���`���0����1�Pd� ����
t~K�_S?Pj�%��9���!�"}�kU�1�0�?��c��j۰ھC�k���^֫�+^v��p�Ū�J+����|{gb�|�P.8ܹ����7�3��IL��@��p�@�xV�2��Z���-gɶ!Q�ᅝEn/��4�/ϴ��=����*8�e�$M^^��b��4��qz��/�<s嗺�J�.@�sZ���
��c��������/���X�@e�zH���oZA�[����I[]�
Y&�8j�����f�mq ����ئ�J�wex11R��p�t{�p���y�^x�4��1, �i)�HKu�7��d0��]�2:H9��<�<F��_NԱ$��-�ܩnÛ�i�PW�����UG<�ŊY�#�w�X�]䒳�$��>X>�2�Ж�v�_�]�{V�J_�2���)1u��7�_��t��&dk�(N\^H�/K�CHbLY�����w���IA؎8�K=�-����(�O���6y6X\�=X�V6�5��>�>����Erm|L��2�?��%Z���_��hZ�ZH��u�������x>�%�ۍ��̎�KD�С�l	�?����0�g�7=���t�e�y�@m?\2�P�޽.z�.6G?W�¬�*��Pb�R�DXʹ�C2�%�-!my3X���}镦�:v���~(Iƶ��R���[�n\e5L�E������,!���ȕ��vv��s�tc	O�Z�Dt�6�	�Ҳwh�k�q<�\4��2X��F)���u�[nk�˹�$�݆���\.*�v�� r���C���� 5P$U�p��?^m�]o�������Y8�He����v������{!�.5u��3wk�2$<��s�8��z���`M�DND��9��^}���N�g[�e�$��AF��θ �n���âh�$�o��NQ�l�:X��$a�a��6x=|K��Џ���"�,_�q�j���88�ϥ��Z��f�z�lM��;8����1�o������~��,/�X���!2+R�{6Vꩮ�Z�lO�jZћ���ӹ\v��_JE��P<��ڏ�X�B��zTA�xi�B�T���n�rP�؅]%W���Z�x���5ԁXZ��	@$$��P�tj/C�u�۰.b�xtz�uX;��l���Gq3si~ݲߔjiE(��uX&H���{.Y\?�����]�݆I�3��.���}#<�P��L��}L��Galf�ɓ	Xx���s�T=�9��e��c�:�Ef쮕�L�c��e���%�̖��D��� @)��7�����Z�2��f�en��*�5z�����`�Q�j���N�輳u�����6���֜R7�v�
�����ʏ�g|�4��2wM`�9>"W}Æ���OP���O�ku����fr޽th����O�Z��땭ņ�V4�t*�t8a��߀��j��(8�x�OA�m<w���I����ȱ�� ��"� )������G�ե���ͱ����u�Ҝ���}�Nkg����TS
V\���o���g� A���Q���y��ﭝ�W^��n��n�(M�r [&H���Á^���#��>��ȩ/�_X~V��m�<쌭$��I����/N����o/���z�m�м��Ͷ��u0�ҋ�eߡ(�3B�fZ�k���l�Kzb��G��3�/��K{���_�3<�{��$L�{�r���_��M�����g���J��?m�Y�h^�}�aQ���ep�y�u�x�m�dM<&�yig�7��no/��\;���6x�u�-�%��Y���ୀW��N��k^-Zy
]����e�Z�T�XEx��S���Qv���l`iɿ�K����"�|t.�ZX/)�y�5x�#��߮\>��_=⽭[@��،�7��Bu����|D���ѭ��@gҜxާ�Oͦ��)��B��pTRU�7-��Rf�i�(��V
��%��«�dچVȫ����G�&��Md{�2]������0�����ZM���gP�ڨQpڔ����J�?��Ү}�.4_����緷[~��~ E���̅�E��0F�R�=����;�%	�*A�WF�����<8�Rx}G��GCț�u9>�m�dI(JR���q��D뺿q��~Z�ah�b�h[�6׼���+!j�Vt4��.�[ces��4��u��;����z�68�gd���9W�Zwjt�/z)H017�M��R�^f��TGS-���Z��1�E�d'^�uwS8�gm����H�r�?M�7j��yū�۝6'8��L���YM�H���6�c�q�C�C�����h�lȱ3�����%�HyP�e��|��G�qƈɦ�Y��Hw��	���]8l:H$[���m�����-@�/���g��P����NUly0s��R�k��LǤr����m���m[-<Bz�Z��0"�s��b�*��(��L�{�|}D@K�-�\䓿`i��VE��E��MK[߮�_� �V�`h�77}퀰�9��˜ks���ǳ�7n¯��ξ�:ףЃ��%g�� 9�t�Ш�:XU[[S%.	*:J�'ƇHߺ�O^M�
�<�|{KtiM�"��s�������q�6ljD)U�KDـ��Q��{�@�deO9gR��]���8�����K�񽮲��ҴC�Vv�t᫿h�s0Ȃx54�B,'Xs�~���-�͒F���i%GV�f���R3ߵ�A�9�L1�:b4�t��V�]�5�����/��U���zřy����5�#��w=�C]��^�;�b%a��4��N���eoC���g��O �2��r2�1��:*q����'kѷ����8Lzt�/*�Ȱ�s5jd�� ܰ�jWC˼v��֬���y��d�9:F��m�<LE� ��t��|r�o*�k�7X�e(�՗F�J�uG�ks���������Ǯ2�mr=�����f#3E|�;1V̺�SsF��ߋ�1��v��Y���z��d�c����uE�s];W��!p�ю��j8~���rF;a�a�n��E}���������g�sp�g༷6�D��;���Uѳ����3�����]Kg�-]�ʣ͚S���~d� D'P��3��)_���	�?�
�>����k�_�kt�*a[�ms���.ȁ����2�����v�2�#�o�h�M�5�?�W��Â�=�-p�U�w�)xQ#}��z�@�c#���'��_/%��m�t�i��́�����~�J�-hV�<��-"%���K�Y v���yɪ���mUg
���������󗪞�-qS+��Vr����ߞ�Ws��	L��J��۵�̄F/�o�Ǟ� :#yzi~!M����(`7S�_�k,������X0�	�Q�j��¶+cD��x䖗�֯5�2��i~�p?�����'���`Ղ��@���޵�`�b��ŏJ�X��#	7����/B�m���\�9�{�ڑ��DO%�����_Y{L66������MV�<�����3ؠǨÁ��|�ڧM׺��ML�O�i�O1�x�E�9��ou>֓�tM4Nq�uAT4�nC���r�5g��,'e;��Ӈww��(�,��K����T��'��&.%i�ݵ��(��^�PGf�a���	U�f��9�ˤ�Ն������� .��iҗ�8�s;��q����iϪ)x�6gO=FU�Ww�f�&a��^�*R6|��Q�������1��k��a�[F���֬"���X:�`�c̳����i�x;�k�K8�@���&:�:|��!`�]BN����*�{?���W�������WR┼w _dO ɕ�퉋憪Azl�����R���Ӣ��Ɛ�狖�P��͸� �p��_[:����_K>�fSm��F�o��q�f��)u-�� ��;f~�ؚ�Ϯ�l�'������ߗ%`xiV��q��b�jR'k5�}3HY�}�5ś*�n� ���?���u[C�R�G��0�8������6��q�2�a�~�	`8Gwg� Wj�z��q�,r#B4	��?f�i�6��>UGS����=@�����W�ZS�����c;P}ѩ{���q�t���Q�����`�ڰa|#<l�+��n�
/v�N�E%6�vl��{^�o�� K�W6θ�����rL���S��8U�����f7�4���b眻LT?��J�W�K�^�	�����`A���"w �+aR*�g�Őj�x�]u�����|�n�����VZ:�[\%M(��(�W��é�@��7�z�`�����F�γ�ra�F�Ix�qk�α3z�b��=W���h:�&03�������4c��" �s t�!�_5x��cC�����]����ĲhU�(e�_�8?�:A͢��Z=��!{���罸Vu��8ƭ*(����޷��6ZDɂ��⍍}��L�����B�c��a���o�r;f����iX#7z5���R�a5���VZ��g��
J��?]�HS�d������!��>�ͶK�\a��w��G-�j~6����_�6�?�QS2��1vɇ��ߡ�եڷ+�8�婇�W��h����J�\D9t��'�D�$b~������Tc�(�
u����k籜|{�M'Wtp��Ob#� x�9�f�D�׏�>*ng��gs%�gw
�?�o<�_7�@���d�n��y�O�o�F3��(fU0{��~󰦎� �uZ�B�O�����\r (���ds<h�M�*4q/eײ��{�a�í�	��&ݔ�=�5*�uq�����
���\��`EI+˷�7;O �藊���1�z�;��WV��-Nt�ޟ����Ԍ�-UEŅ�V�La���8�@
RU�yH��� 6��Y�3珮<8Ȱ�Hs��ד�k�E�m>�1C��������BV�I���C�qx	[{F��f?WbF�Í��	�v���jS�(q!W����d(%c�`b���-yOH`ٽ�w?J���=�3�6o���h�#ضP���z;Q�;ߪ��n�~g��~7�P")"՗X�����m�l��~�����0��b�"�o�Lw�n��{><�	����C�y}�#?g�-����;k��AyF� ���c~�ԖC*V����k��me`��r���5R�gf
�Nh���O�f��%4`�Mn�. .Ļ��mU��'��
���e؍��U4�z�!�W'�#����]��ƅ����C��e^���>6(��q��9�$%Q	�K�4� V/����qhG�[�)c��YB�zJ��qn�Q����1�k?rp>n̝��}H&%io��UfǗj ��w��Z�8����čӂՋP9W�๩��&�Gs���ٞ|5oɖu��\�^�٨�f���r�;�ct��]I�]?��pNJZ�G��'�T�Y<B����aĺ�a�߰4^v �Nj �m��~-[=����KB���QS�2tIlz�WgO(�ݔ���5xi�d����B�?��T��_!��;vbC��F��+���K;[wh�9;��b����\kۮ�x��9�ww��-�H3m��]���r���?��>C��S?���B?+��0v�.�Үr#����*�9g���eY\��A�0 _(�E���|H�ۄ���%Fm�I��ܮߚf-f��oo8����X5�{4�����K�+�I�	��mvx���G����o�a͠��?=���$A\�k��,�
4}�����6��f�f�X����B⫝����"�UxhH�XuyY��D�U�-'�L�P�O���ݞ?O�wێ�['�\�<{xs�4��r��#Cv^�{�,�˹߽�X����қPC���F�\�n��:t���_���=ks�7t�QJ�7Io�hb�S��u�pX!qRE�*Oĳ�.�6;�#���]�lV�{Q���NG�:mJf�$�ѓ7��Z|p���̷���W�"�������[��t��t�&�l-Ky�S<��a�|��iJ��qK4�BB��iɗ�xU�n����#m~0q ����x��a�)*�N�`R�?���\|Մ|w���I�Ms_��"���	e��i��Q2q y��JԀ�M_��m>��e�f��o�i�T���R��X#;2�De5�_�j�� ��a�6����~b>=�Ԏk��r%�-)�J3��zl[*�@���.��D4�[/B?�*��}��������<�{ػ}O[`��e��c��&r�Q�'�y{/;�W���"���*+_�4�:̭���ّ�<E�1�o���̕�5y~�
6V�������?H�~E������;�c���ߙ*8{],�Hi���*�5h?�/}c��䯌ّI��ICy����@O C�z���T� ���g׼͗e��7C�::o�ϟ��u��~m9g�R���%a��KgK;JV<�O�h_Y���?�.���&�<�
�8�}0��`<����9��{���D�n�	����$W�}�t����&�d�@e�K��$���p5�U��/��FM��8��"�K!lB&�OG�M�>:d��Fg�OFP�7�a�<8�N�LNG��p+_�]uE���q��U�Ц���$VdD��}y�k�K4�M�,�|�t�e��\�A�@�!�'���&>��9��U�����~߱��v�֯���d����线c�7�L䊮	��� ��s�J��TmĊ���\��a�D�ӊ���.6�&8�0ߚS�=j@�ʲI�u��E��.��zIcvox�b����'�'���F�GR"��]����z=��GM��(t��<M(k|Y� ��?<3� Br����K��h�����MZ߻|P6�A�^����&��0Xkz�Q�g�4j,���Q4��1���8�������U�Z��>��<�0�
�,B]�����[����9���Ks)��/�h	Im���	�u��W�ڑg OK��X��Q���'�g`��
�sL���'����v�9#Yq����:b:���	��&F~P��U�3�85�b�P�_���?�O��P�j��{�t�����v#�Ņ�"b~^J��A+�6��Mxd��L�;�)�*�ڑ^�R��?e{���nk����c0��4�B�*�vM��x����E葊�J���'�r�Wz���1�2�1C����,�<V������#����Ux?u��N��T�G��/	i�"��c�f�Yj�,�;�[�aϭ�Z|Q8�q]��˙����8MÐc*q~6��qͽ�V�IGǾM*^}kU\]d4SA�;����	1٥jG �t�� � �./��o<D�*I�p����4��[cר�T�!��6��e��_�wġ�?8󆴧��C�$`3I����Ǯ�_|����:
Nu�qܭ.4��e�@�h����'~b��� ~,5�o}�c*�+�_�H=�����o�ô�2R*-9�ҳ�����.{�:��j~:рٚ�v-����&�!P�9+o�ql�j��sq���`�/���۷]�� x9r�Z8�$4m���'V�o4�$"��B=M�LۺѶ�Ѕ7��\w[�s���L3�Q&5q��%���/���Jo�s���N ��7���P����P�t��o?��c���(���E�W;��O��,:R���Զ��>x��}���'�`�/44>��%D��Ϳ����mN��n�aB�=1��)i$��\I�#T�����sx�C���ks^�k�7��m1@�ߥ�U��2���+h����we�e�΄]�-��8/��.tKXM�8��c�)�O̘��ĸϬC�%a�~�̟�Sq{�"k�钥{����pVJ�W����p�!��s��w���gԑݯ�9������*;�،-�-Jd�G��ς�Y����qw*����=�CJ%�d���q���ʹ����E{P~M��+�<����%�W�����}��X�J�[K��!>�"���L�)^�s�ѥ^�H�tk$MU�].$�pj7V�-��H<�'j;K��h��� �	p��:�%�%�w���J�TN�����wj��\��wߪs.7^�Ăn��������j2�:P'�G�\�AV�0�Ȼ񫔞c���rޠ���j��u�!�B���?�����x#�1yC�g��Q9�����t�N?A��^5Y�Dq��/�=M��e�ȭX��mm�������Z��{��h{�qC��FbV�dvH�v��,�4���X��bV@�l̳��x�t�^�?Q��V���Neg@��l"�|�p�k^e��l�|���o�~pO�|���9��ˑ���%෸E
{�""�S��j�ѓ�wm76Ǟ��ٟ�g��˂�����؛k�����-�	�[:���E�#�w����w�S���&V��ݶD�C��XE��k�0�(̶��_��xyM;�5������4q��S�	 O6ܒ�,��!�P]	3�kW�]&�����ٔ9�^�;!����B�A�el��[��~�,����<�±=�~H�w�s�zS�s��c�*�lM���k��Jp�waCi��cx>�k�+�6!��ب�P����%J�u��3�Aӥ�j�����&Us~��*R~�"�I2���+s_{?���Z��z�n<=0�����/Aʓ(�,�y���sIq�}�=U}��M�$�VID�@ ?FH�[�If)��Kj�F�-S�tw��q+�-���FN��O$�%;��5A�aGH�yƲ�X~y����-T��}OZD�U�hD���� �/�)��d�H�5�qy����ǎ�ZyGFrQKn[9�&�_�Lh�RXBQ�����; @��z�S��z�zI��初ɴ��	�9C[�r'�߷���k�?#+�_ ��^�ڟk*����7���[q ԽŘ�R�%z�Ml��5y<�x��KW��󹑽5a9��M#���"N�ɀ{��<4���?�`��PՋ	M��O�\��������1N`}/��͢7��s9M�>Y��G�BYj�^iӗ<�']�h�I�_��ok�hv��	��%(|����o6�'8<v�-+�uZ�}����B2�li&���v��3w��RfX�E������e���9o0=z��VU�����e�kd���\P=�V��
�݄�D^l�r�ud��&�U�Ұu��|er1�P3ٕ+��aμwu�\d�ⱠN8����C�T�7�3��� ҟ�'��=�_�k��<!QO�ѤJqOSˬ�]�^���#�	�3�6mW�\Q�ڥ��g`�D?���)��z�Xq KB��|�z�s���px��b���Ϳ�����x0\v܉ߓ̢>����'�n+�����-�ӌkWd�O�u�W��v~_�z�A���ڝ��sL���a<b	��8�����ޞxɓ�3�-M¯o�>z�����5a�����%]��&=x<��.����	�C7M����"�.�a�4ƌ��Tt���߫����e`Xt/�W�'A�Kc}e���Ufŭ�ogb�|b�1��F@@���e9b!,��&��_kqPx?\Gi�F�:7�T���rh$�o�Ҵ_��H
����LJ�����5y����\���Q58i,0*@���0{��3lg^^n8F�,�WGLmkuNS.!���9�Kzl�F"K�,7d�/�e6&om{�{��#ʿ]_�~�釣²��*�K֌cק�k���Q
n(���_���,���Pɸ���q�Yt���֌ğ/�R�1%�*�
�-��8�Í�a_�Y��RTbM�h+���\oww�6K�cX��L��5���1��1�֥g�ߟf+���]�'��:�;OH�]�W�۟����}WX�[n;[���m�^ݸ!B J(�0D:���*-J� ��B�(U!�P�C�-� G���s{���r�'Ϛ5����7_ր�Y��S
�*��jUR'-���E�Һ:,�F���b>���)�TU�w��֭�`w]�H\*hm/3=�>>s�S�V�1`��@|�����Pb+�*����=j~n]4��w�'��>QF�7��0=���G�2?@2�G��Cnw��z��&�p����S�av(��mXNfN n�2�������v�|��GR�;����@�p�J���YC��Dpa�}��/�D5��a�|�es�b�u���qa���!�?�5i)&4SV��t�('��P��l������ԇ9R�.�9^f��sF��%�p�`{��vZ�n}भ�ې����b��\�%����P,8wG��K�=� �;;�!}�V�E�?�㻃�/g֮	"7O^a�>���{R���Y-��)M�z4��.�쾥3SoR��z�}���n��h�U��%����ru����3���Ǔ�F��h�X<r�M�� S��f�=�p�+��2�˂�B#�γ�a�7ϗ��f
��x�|��m����}�3����8��O����k��zg��Z��λ$�9p"��՟e�_�L��tc/V�|�T�Q�ԝl�_A����냀��RIn6��<��S"���C��p�W�C�����1`4|��|_��'&���r�f�_hӶ	��c���p �%�حs�F�yǌbĵ�]8�7��mY��#��&"󨵗�,��]N9��f��Mh���us���q����L�[of������b����K(�s٘X����5�,���8�A��5>��4��V�*7��\�Eµ5zU�!�q]u�~����9�8*�,����/ަ,��;���-�Do�b�̫�Y�}�_ �W�Y�2yb,}a�!'��ɼQ��t~����K�)��H[�Two�t�@HH�H�H]?���E��|��,�1��vB�K��&;K3#]�c���dxeJ�k�[v���v��T�'��:T;�9r���B\A��`���6lU�?����H(��py�;��,�Y�\A�I�B@P��4�Ű�('�;ɖ��|0�6���(�����gYϹعW����	ƺ��M�\{!G��8%��7-!��;]dcO���>zݠ����7�76�Y�ŗ����?�T��Vs�<q��Q^U���&Ms��F��*&����@a}�6�����r�?��	]��o��<�9U�XU�ك���<<�j��Վ����v2Ǘ��.!ݷ+H��ul V���|&�j#dbJ��gC@B?mIk?V���c�ʽS�hH���7 �_ȱƚ��jO虳ݺ3�cE�6s��iq�D\~�%#F�׹��k�sz,���`���)�U���Jn��2�1�YdS�m"�Vn}S�{��ڨyԝ�9�P�������<�(S88�W�v'�����q '��1�T�IF&�fj��� ���iV���#3���ǀ�p��M5�����"xM���v��k��"�F�	y�<Ý�R�(q+ PEC����IRd��̅$�t&o�Ҵw:gmEd�k�`�������l��g̨
+B���4z�`]���Y���	�q�`�J��w��VU͉֯$	m��K�F G���4�vw��Bo�E��$�#M�<ds�/G�|ޠ�L�C���CM�'���xs��XI��}`����kIT��E0V�]��Ф��a�_��E.��d�a2~T��K$9�]��)���.w���)~55��$�eN@�ϱ`яE0��g^�6�?	�)��R[�ͷ�·T��y���H������{!E�����9g,^dpA�kae���6
���
�'^�p����zXO�^���%-���k�x0,7[O��|A��H(�o/jK�� .���e���~<��y�Ts�3��AJ�C����m��R���Lm�<�Q��EGĽ�=]ǭ�2��H梨w�d`-���w�,�K\��맃�e��(�ٍ�D(�$Oh]7.l��-��E�lȶ7�D"ֵ���W�{߶�`vf���_{u�)1*^��4 '��$����P�tH�_FT\苐�̂oM�H�*_�m���g��Ś��\���l������*���Z�~��=�z&�:<�]pe���eD�Qb�=^��潀I�D���/�(�q�� ���/I�<�(��	��q~��@�W�;�~k�?�@�%�ݯ��^vϰ=�$k��3��XF�����p�}QӠ���JQz�6H�
�]7�~�B�_�����-x����ȏ�>0��᥵7	٢1�%���|�q`�ܻk��L�@z�&D���Ms�~��2��ݜ�gf�b>�,["\��?R���^�Z�V*yH5�<��Tc�qf���(ݛ�l����o�9h8�� 7�<��vr�Zh�'ō�5�;j�e�[��sh/�R
X����F>*_�e���]��T����3�������m1H��L����㦞�e�FcƍSG�R�qT��S�|�Tϣf+
>/U�gn���{��d^�76� �Z�ʬ�2u���1�6�f�t��~���q�6G���L�[�n��~$�N<���F?	�V��L**�1��Q��;��4�4�]z�s���ͻ�߄J_�����pCHXhv��M�DTbֲp�gy�<U��0���i�tI���n����8���'�������aN�V�6�&It��t�C�_h4�r1u5TJӎ{6�J��m鑐Ƙf4�42	a*f[���D���>��(����{�Mv��S2�n�'W/�;�R�qtL��-�!�rS���s6)�)$��n�c���Xza,t�����'��������%�k��l�˫8m��k�u�=�`���:^��Z�ڟ
n��t��m�	���V��u٦Nc�l�A��"�������f��|�[�	���}�|��!�vU�n��b��a���m(u�K�#�$��Ҧ�,/���4�PoC���������x�\�~�南��-M�Z`O:�Ў��.����������~w��~pI1�f{����~�w:�b%'1�¥Q��9#3}_2�cwgB�}+����ML3�dqe݌��y�>�&����nPU�_.����i�ę�&��郼�'�`��?�;O�*��WO[ �,��L�iS�7��=r���E���!(>�Ӗ)�'��O.鬆ϓybM��זULLg":/�x�|h���&֪����,�N��(5R��n�4�4�$3c'ÐS�L��;җ���)���e��|j3�/,�Le�D!5�Iy�<�1�͊ס�����9A��>1'��#x�˦"�����H�m��@�������T,�Y�����H%��o�t�������\��q~j�ǀ>?�*���d�2����s� 	n��,J�`�D.x����t��_}�̊o�TV`!/���9�^�1�?�Z7~D���8�C�ֽ�yn��}bw�37��V}Fx�����xD_�����剥�Ë���iqa"��6?�����=�]ɴ��٤��W.Q����[W�ʆ7W�v�E�~B�w�%"z"��~��f؎^d�nۨ?�B���^Z8X���Kg��@�vY�w�6�h�f��wn�~�I7�y�挏��O� u3�g&k�(��)�6M�$a)��t�R�lR�42�yw�����ѹ⚁���J�)!��V��6 �cΞ��ț o��h���y����^CT<^��$O,�4Ó�K<N@�;��CG_�֥c/T�[���1�s��D�H��F�0W�B>�l��t�>��X���/L���n���p�Ti�(�K���c��ؙ�B!�
��8��'d��QiOP��>3���ci�׿�]^\Nl�4�'��Q�����%a,皹:�9��5�AW:|T��gm�ܭ!�p�f���n��f��J�P#-V�Ǹs�n�ȍgtup�����V@�.Rך��QS^�4 IB"�|��lw�;:)��n������k���ѣ�{)fD�n�w����R����UA	��+�{`bE9ܗ�^Gyx�%�W�3.��d��L���T�m}���J�vS[�S=�xKyd����{+dx׆6t{�����|9��Zɑ!��/jh�{��s���������,�4REe�4�nv0�m+0�ͩ��kn=�0g]4[��@l�s?���@!n�atU���bT�{�����yK����]!�1p`�!(3�A�>�X�����B/���}�APWѨ����DC�X�R�U��=�K����3;i�XP��ImY8���y:"�4�ASTL�{�,�78��ǟ��13Wc%=;F�/��[�*�ޔeЂL���c�^�[��B��ƾ�J���H"X��)f���ґ��sp6��`��ky�ۡ��CqS��*�\0sL�ж%�F١���v�ѪQ��.�)�5�^��|�÷�'�u�C-~d{�v�Ax�/�z�(T�����v+w/�@ #��@�@y~-T�{8�b��1�2�6䚼<:�ҬWg͈����4+�+�ps�Σ �%�K�ĦY(�c׆�Ze�,�v���	�F�΍�3^�Y�#ap�<��1 �T0oO�I��R�*d�S�^~��'>��۩�my ��=��{�3�$����;����\=�?Z�Mɩ�c�Q�+A9���V�%�\�"X�eN$|���|��LU�A.I��S��SV��Z~Z_b�����w[>)�g�5�P;2c_|/qq�I���aBF����%�9��I�럖	��j;��%j�*��-��~Y"���~����;�*�����V�N�V���L����RN��㗤�AJI։|n��l�2�����C��f񧖸��o/�[h{��8���"�_"�SR>x�c2�K���`ˤ��(���G�Z�}��HYMU6E�s��q?����h~g �l�T�>}=yi���>ZiV,d(�XBvS'r,���j��*��x:y,e?v֪�z���ߕْ���� e������M#^��M0�������f�|j7��@[E!�TW��=<�}H0Y�2��B�=���A�8���M���L�wߗ�;�X��a�H�T߯ϵ�{�|�!�s� Ie����\�TJ�o���]W3m�,/ 9�����g"h(����TǙ ?�Ռ��I���ď�Ԅ��W���moIݙ�N��eg��&�5˧u\��iӷ�W��,Y`��'��Lޥ.hF���?��z�+�ԝ�1vۧK[��C��r��,����&~[�|^��SV���Ίo%+�(��׵	%�E�>��ԬMA��x���Z~� {W���Th�,�q����C!^��W��$r��ܚ=�1@��dmY��Qf�[v�̻�@v}`ߓ�'8���P�媈�p��� uyz|]����m�OҮxm�1��F�K�:�+���g��$_.}���R_a�h�y*�¤�
��%'"�F�|Ot�9}���{����&0Ӭ)����K���%$��T���|�|:}�k�+����,2!n.���(�a�ciͧ�k> �%x@'��3.��dvQ9G�I2��Z�km��I7o1_?�J/���tԓN-
ys0���ks��9����b~
�8C#R���5���8����
M�q�4���
�j�� ��WVRW�H�,��4�:z4�Q��	�H?�jZ��x�a����P8�sҴ@R�{/��;D���YQTfL׿~ޫ�}��(E������n���W�<]g5{�eU�3'����%'��mi2����s���>���m��^����:�_��[������K� ��5AfɅU��/�{T�5�����#y+��/J�y�h��KAʯ�������{/�z�{��\�����Z~(`%=����ӹ;���j,�QYB��M_���3:��N8����KW�j�	����!�+epI�b5���8(1���
�0ڈ��f���Gp,%�g�"�M�����C6�L�h�u"��HȻ�`~�@.�;�u2�1�{�r�mgց�h:�n�>זXwN������]���E�����#��k�ǀ`�*�QF�m�#��n3Ni8
J�w��}�7*�M�':��MZ!T�v��xG���0���(��6@���56T�
�r�s̸ٓPY�]���N�US�q�DpS��/��� 񅒭����(1}1�ދ��Pk�NeB��1���2�5�fQS�_g���ͬ"?9UY������Z����h&-�9,?@i�(�nVWd#u��f��1�y�Äz��2q��$~�s�S��3!8�����G4��i�c��,,�+��0��q	|�m�ѡ�27�>w�-q��oVW�k��WCҀ���{/�y�8Ō����Q<��60R�h�iY�σu��ʵ>P��n���{6�=�<X�4Uxȏ�n"���qa�(�=hڳ�f5`f���RR�dޥ� �$[5�?/"N��6��ׂ��9�=eъ�/;$��|IvA���m���m-۞�JT��������#�ci���bkYÆ1���P�3A��x-�A��A�bxYd၍�Kd��-�z���.`�P���W�Y���W�~����{�����-F��5��=Üq������4�[FӰ5ح[|Ch���y��gh���KXoz�}��x�~�c=�\��*�Ki�CGc���g�rhu��J�hJ����AB|g�Y?��w��x��`�ukZ֧�-YNk�螠���5��&jK[A���Jv�nt���%O�k�̖S?��%�d�/�774��R_����ћ��Ǹo�}�QgD4�nL����0)e͍>��L.�X��:I�n���Aͽ�#wu�*�I�UN'�=2�I2��k�����%BD�z���r�Ւ\�����@��n���کI��~��|�/�o�*�P0�~Ŕq��&��B�N�o��n%n�R,���:��&z4�Zn������t^��֖�ʅ��Z<H�n���.�2b5Љ`@N��7[=���D���N�W�������Ǡ��l��#j�	V�㥃+cw\A=�^Wƻuyū�>W�,�`�`X$y�I�a����{<=���Vsz�R�'{����bH�Nϱ�Jiw$j)=��v�|����X�]cu�a��ʄ#?�ᕨ��S�թط��:��]��V�)��&S�w����#����"�]H�,+��_�$���4�%�y!0?�ؕ����~�i�^U궫Z'��]ٻ�b���`�"H p���8�{���L	�/���!s���݇Q?�!/������gxp���:��o���y0���b�G���*Ma�ԃ
	�K3R����cf|Č���T|���Q@�H��I4�c����4������z���b��~��K����f���sJ1����@:����VifEf��y�e|���ܯ�EW95�v�b-:c�ۿ�)Q�9C[���u�������fQ��C �b<�%��O(�,9u�eo&�g`�UN\⭳v1�UMR�	
�3h����G�J���A+_�(��b�8���z����~*\XđTX�E���/�*<���nc�t�?E���2I��N���g��TN�ޚBR#7�>����z�W>o^�u �ǒ�������%�J���-�ȾFW�Dni��~��dL��ClMe����O��c���l}�>F�ۛ,���r�C#׬Lp|���� ���fpL��̫�v�w-��O�?��$p��R�b!N�q�@�[�=����?xC�=�W�T?.��ڰi[*��8����H���
���f=��"7=s�mV�H���������/`��7��;r3��2��c�8ԛ�.�Wl'e #*��omjAL��J�"[�潋���L��4ԭ���m������w"]f��eIj;)0��	�{�h������ϔ�>�(.�@���R\m�ab����qz`}��/�����([m�1�+7��*kt�:a�X���M�K��D/����<ip�%ݹ�d����H-MA?�z�e���+!:nh�!a����c����m���-ca
��j�|���V��v�Zm��Fa���=�덞�Gv����}+��E�D�W�����	�Ҙn�;�_pEnU!�B6�epĐ��VۖtVgs�QaV�=�Гn����&��U҈9
>���պ���EF+����%�-4������CR܌��T��ԨG�����n�lջ���M�wk�6T�t�(��*zz����
����ќ��1�:��Q����k�1����(3�U§˫vZ���3������6h���[�m��VN+Yv=>J�7��I�x�Z�`8j-�*�A���U.k��TJ�td��<�xx��?1��(ý�Ų;�l�)�	�j�t�>�����ǀ�������MT(�{ե�	�*㸝�U�����K6�����R
�f��棋���J׾1b��BB��|p-Eo��� o�Yչ�	4'F��e~��		�ﭜN.���Җm���;'��m'-���h��<�$E����)e����A	W�>슎:-�z4|S���@�N��P��.Ȩ,ڇb�������ʤ|��Qo72U����'p��j�>ݳ�iW�M�#��0`�A<䈞�
�-r�������Ŷʆ�NnZq$훑W�+�W��Sy5"���[b�"-t�����$�󫰻k�k���1K��;D�aϔ{q^�m��Xu���!0>!8��' ��)��]�(UJxIY��W�qr1�� �^9�����|��A)�ȱ(ܳ.>���5��4@������(=�y���P5żO�e�l^^7��j�,P�D�VS��f����a_��~I@����Unvԋ�޶�X��WP�s)���%ֿ'�؆�9��t9�ks�;���Xh| N<��+%���C�B$�\�o�u+06D������若�1�yG�R	H��Z5on?YΌ�UPki��������]�d١:��+B1����R��jV�ѳ1���Y�-��;�����sr��t˃���^~����|�a����G¿H
�o�r��^�� V���@�ωs�ʧ��K t2�W��-&(�7Ō�'���#m�q�����M^�RC�5����\����B%�>�F�>uޮ����~Tn7P�~�&oI��xܑsx7��Ҙ-oJ�4�Wx�KR��T����+Ő�u4wW���?x:o�E禘e3ە���-T�/��-��aC�vL�v�k��x;�2��s,�̹!:b(ҫRk�uax�7�j��6��]s��`��ܬ�1Po�zv���(O�`�)��z&K���hՊ�VG�D��6s���J���
��ͪ���ھ?3�JT雝SL��Z��׆��_��'�)���Jw�{Zx�M��X��W>n
i������D����N�ؤ/��fh���I`	���e�H��F�W�9i�{a���ѝ)�{���<sD�ҪL�l�:g�>NE�Erbk��k�!�b�4��S���޶+�%�����P���an�	K;G��5�$�WZ���7U�b�����|^s+���.CX�,��l�%H眞t~�j��sɮ�3ŧ�*�w�yM�����=�2��mG&�H?\��[��ޯq>���do���c��@�s-����imq��4��G�8r�)Xך�̮��i��U���P� ��;DE��_�Q�d�fd��l��=x�K�m#�5_�4��!��Lz�tO�5����o��4g�($܏/��n]��oó��'��u�A�1@����qH\�l��~We%��
�c�)jQϱ"��1OGL��6%O�KyI���g{�(� ��9�L�3�9l3��m�ysq�~�����)v)�P�ݠ�z�(� �P�q� =��˹��g8�Yi�����$m$9��-NH_�k`r���3HD:.~�
1�P��4[辌
�a�0�� �����p5�to����>.��q	O�_Y�I���(���x�^��Wԩ�@��LX���8u�[�	F�!~:F�����G)Y��d�@
z�	45����g��~os��O��&n�w��I��ޒmm�����)LgV�����'5�s�笿`�i�H���_��|JEK��'�#�(a>Z�1@!���6+^4$���d��U:j��NQU�0~���~y���ܜ����cI2i�"����=��3|�샡���5��j����G`�LȤU(�?=�Sc�����7\���&��jɐ���͹��'A/3��󜎺�[8W���
5��24ن���j���}��bG���u�A�W��i)ߛޭ�=��}�#^A�򖲇�W)� �����1��k�ߔ4�;���JZ=}V�鳊�{�t��b��е"�L�Ư�t�y���k�Rt�p\&�0�'�������;I�ymz�Kg�'9-LqZ@���<�G����u�i�}�$e�^uɲ�����T�1�y�r+HiS�A;��ŷ�G{E�,S��gL����X笓zϺO�A�G{T��4۴�����[��=����9Fl�w6�E��}��l���or���}�mu����������љ�:��D�����Lġ%�����"/_��kSu�tN|�ՠ{m�W�Mg�g�`�*"s&�gh����1i��b�֗j��;_*tO�j�Q�D���nX5�Z9�"��E�@��bY�^����{������De�Ĥ-��[n�֥J���-u ����FQfV�A�TM�5��b��)~7 T_k��R���󀦝�W�ƽqΚl��&�Dk{�P�'t��	��]���RH�aׯ�{���]�٦^b���dx� b�pN%ZT[Y��(��#��������ӯ����mj~TX�-6��T��� $��x�`��pn\L�Ir���Nl�R���Y�����3�"��\G�1��1� �G����q�w���lEJ��l�r���{�k]��A{?W�B��5�,6�Ê>V�+;߶��ǈ�Ż3�k�j�c`Xv8����EQ+si�_w�@��!�_�< `���V)�.��n�h׿�`�jL��z�Q%�.���bY�,f���F�aZ�t6��jS���ܸn���u���᝛��{���X�1���~7���mLJ�TT$$�5�����7����F��Q��D�>!��a����9D/�K��H�X|:�]Q̹��WȰ�n��bBQ���#���6\��p����h7</�����e����u�&�T��F�	�V�t\47GJ���ebR��4��N**�.p��nD̝��xH���Vn�Z��|�r6��ʪ�x�w[q�2��Ѥ�Ӹnw~:�sc�$bQ��^ j���m��V����:0�^��z��B�п[_�Q�/\J���<�L�)p��՘Y�ˌ[S{B�mׁq��,��!���&����.3�]���d9�I�߲�/��.��PL\eH��^'<��|�y����\E��!A�_e/����	� [�UAn]R�P����}5���_���u!"^ذ)]U����Ӗΰ-��G�:��3���O��U��>�Z�+�jǶu˦��v;׶�t>��'�7�k�F�����X^/��x���Kb�� C�Pl�BD�!�k�U�M������nZ��b]T 9����,��S�[����$�G7��ѿuTqA�7�߂�,@(Z�AP��|"��xE��ھ���*h�]���g����xd�A�ppk���*���^�Z�j�ׁݤ0�QOEȀ\�0��,*�+0�0EԒ�[~)>ǭ/1�т�j��u~�d�oÊ��.��Q�ڸ$��c�4�ۭ�J�X��=�#�^i�1�Rѫw*�֝k�����s�n>`+��H�
|�^��C|u�j��A�;�s�ʍp�E���r�j�9�B��3��O�i��gJ���D\|�I{��g�qC���O�Y�� }쌅a�_}�o,�(۰o4P�k���i?덼�|=�P��ۣ�k���� ��\�^��<ZK�z��#����gy��G@\��^�PX8�?�po�`9!jr�.��p:�`�����l�}�s8�^�$�h��)M���:����&��c��g��7�L[SXJTR�gA����>�Jsi��(�����Q�I79h�1�U�.�7s���Ë�^G�#��w��.a9�oȄ�����1�&9��#PrZ�0$��.)ϴG��$��s~%���L����:A�~��
��wr�>�U$���
L'���^�z��"���R�8��:S�_�SV��f՜Ji�n�ݖ�D[���=G󥶽���U8��TBT�~�e��mf9�j�~7�^e���l�+�-l��`:Ta.�wJs~`j�\C�W{R��2b��^ԭ9�m]>�#����c�Z��,��+y۾�?�A��	����%#!������B�f�<��9YInL��	BÎ�O��}�ǈ��<Cp0�w^爀��]�~�cD|lI^�_�G��x��l'n��l��
!�@8���x$�	�s��W8e�V�W�=����lu�n:V�G����Dj�Vi}�!�֚L殊/�d���}�\����jh�Jq���H�cI;�&{x���!�7�}M����Tz�b��^T���Ml�ÅVЊ�d���=y�YD�Gؾ����m�}�����EG�_��mJV��>��Lw��Y`M%�b�e��i�c��nJ�<�j�:o�sm3\_9��P0��1�Cz��C�W��̉ݓd(����x�p���
���X�^XQ��Ԃ޸��+���[׎��*�F�e�X����y����/����t�|�5������ׁ�I�ʾ�og,�)����£�q}e�3F��<�h��ҳc��ks(�q$�E�
|�-"Ҿv�z�˲E�eT峔�G���\&O���Z�P_ـR8\���l�J)N���_Q����U1U?H�ͧF�L��Dk>��t��}�-r�����x���5��O�b{��|���=�4��~�lF#W��u�h�_�xI�?�M�p�<8�7k��y��zo�`}�ְ�'Iؐ�t%����%�����p-A�<Xќެ^cӽlə�������p������%x,�LRJqk�����Y~'rgG��Enpt���L93�G�.��K��sP W�w��1��s���m�f�ǟ0x0x��7�C0�����V���q����d�(q��p�.t�������IB�{��VJ(C��1Fͼ.��e�{i�Al������1`��u@,�� J�I%��!e潸SW	'�)7�?n�/e����2����EHtل���kj���*4>����*q���^?�"T_��%�-x��Kǀ����4�DEhٍ����"a�WMQ{���:�W�c�%ξ����Ǹ�U���u~:��R��'D��Q���� �'/���Zg��ȩ�z���n�b�;ֻw��
��K�E?��Y�i�H$�Vg���3$��<T�f]a���z�+�?=[k�(�C�T�c^�ɡ{	����H�m�3�j�ѫ��bI~A�Α�(���%B"�M�"p�5��}O[n�%Q>��v��M�K�����u�؊�qĞ���)~���|2Z������1��#ug������;���hoc�e�Z��t��ۑ�?>��x	��x����d��s x)5$�0�;[֦�ë�Z�����+B?_�hx��&pm���6W�Ī��Ƈz,�	SE?ZK�Q0��~����ʵU�.�8�g�4��`s�pQ2��/i��?<p��)�wc�\�<1'Q5 ��ܗB���!t�V�ވ-�9GT�=
nMп���tE�Y�UrV�^�<t�K�����a����0�+�/Dd�@gs��^w&flA��˶U�)E����ye��!�����_J{�����>[���Jw�SQ뛁l�l�%���=�6�ɻ��=��EE蚯���e�
�G������W��c�z!�h��E�����Ui�%]�(�.�+`�����ے�q�k+���z�P�5�W,Mk���/ݒ;x�QI_�����Y�@��l�#��5yY���6f����O'ϗ��V��t�Kˬ�˽���dD�鎻:�a�Ή���gu���#�b���g����*�Büz����y9��9�q��v�;3���M��<i�ѮtzV��(��Ca�c;�ا�i86z��������i�/�S+s�b����	I�)�)UEr������_2I��&�#��Ӯ�d����~����n���{��*Z+���R=��d�F��W5O��O@|p�QIl!��g&0V�*a_z�d"�����V'���V�wЇ)�*b�zU�aP�]��5F;��|�5�WN��W�܄j��q�6�.�9QD�O| '�xgNd�|�T��x	�E�:�q�+t{t��<��O���sԵϦcs`�U_ܱ��UP��|rjde�%��1m�*2Ї��<�x��b�%'�Ҷ;�,���;�8/��G��V���eTN����C{���
 ��u���@T'��Og�^iGT ��h��B1V�����R��H��TVvH[�M1a>��s�N��[P4g�+5OM"��?ե�ʠ��H��.k�F�Ʒ.q�;��l�𹡁�zq�1��@zI�8�\Jn���~��2�v$c��+���t��i�͕���Rw"�*�a�����ztc�J����r��VJ����!�Ld�|�!��ld�,�s��:���ܣ`�G�)�B��>��9+=���w;U���3
�Ϙ_1j�:��S`#�ӃMp��-�9">զu}�i{�y�ސ������2��I���<~��*\'�Œ9:��L�0�:�Ў[
��Dwh#V�b���^u�v�,N�ob�u7���T�����{'ڃ��by
�A5�4jg��yh6A�{\ݺ'���k����S��W��^f�`_�OV�u=������Zu��]��.�Ii�!cd6N���>��K�xy`�Ea�;�H���t5%�����ƴ�vLȻ'�K0KRb�<��]t#��F�U�49`'����C��Q�I���r�N/�l,��ege�"�f��DbP`29�2���Y
�bE���"f=��������1	X�v������;[��{�t��P��n��E�Y����M�%�HŎ]�@�=k��}�H�+c��Eh�V�����#HN�Z�j@�9��ub����<��b��CtЏ��0��w}��Z&�U0+�ٯ�o���H�Y�ԝ�hk���j53Lf��F�w���N���kaG�rv���	��j3s������<��kf�</"�=�Ւ�!&���["�����ZRKƲ�@tؙ��tf�>}R���Z�5k�W��U�ȌJ����p�k�����>�N�seFR����|w�v�U�%-AC[K�_�kү�o���*�*��-P���E[")
��s�u�m|��T`Ա�M����n�}�R�����q������J	��S���N��iJu�YS4�;�W�*�KQ�+��KS���*%cb�4M��C�s�F�z&17OUk?���MJӧ e|x,Z�"��W��Z�]�c����e`��ܪ53㤷Mh�^���,�d>쵆��E�����Es�}��6@�|%e�>��Z�;q�����>-j�H�7�-���U\�4lWg@S����1p���)��K�o�sVkE�E�֋�9h�������"J+����Zee�G)��U��k���-�p<9�$��,�	;g����7['�H/<5u�&���%SĽ����r����#	[��Z1��(׳l@� �<�}��c`��(�Y4�]r'I*-g�y[Z�ȯM�R��$�
{������0�闞�$7[�h�}�;��3eh�nȪ�nҢe���`�Ӻb����ñ	�����/=�߽n�b\�[{���,�5�z����c�:�}V�Y����9m���~T&je���K͡-pVk�M�?�����������)�ǾU�ƍ��o�%����2�&�k>�3��{0�����9����6�}ګ2��T�l���xm(4~tzo��ztk�H�]vsegBB�x��]��N��m�8�͗�;��1���8���UK*ʶ�g��/p:�2��	ey���X�/-!�x��t �Z1`l����{��������c���>�c�Os؄t�V-g���@R�J$D8���=��N��|!MQ��7�>�
�L_�_H�O��c�ehq�h����蝩�l5_g���'��\�������;���bjm3�5�d����W)e&��)4^o�?j4��)Q)��T���9�J�S����U<���6���s�J4ܓ�Og�v�[B&�ep`rX��r������(��$���f�l�e|�T��������!���H����p�aL⃤$�
a(��+�".�T��F�=|5�����r/��UOio}�6b_�r0s��,��n7v��Q/�	���9��<�S�Vӆ�iV���}m�����*
:��CD��^ؔ�jj��b�e���c&����>�Z��e��*�Ǐq�m���s�g�g^~���������iU�uTC�S�a�"�y����Z��o�8�*]�v����j����N������AO�G�U��"��]��(`��3*�+��^}4W�c4�����噷Mt�a����:4��/K$�v*!�`!ՉK�ޔ�N��.R{���.�^9�ֹ�2a�r����b����ph�]�}`E�����?a�~�_�CB��D��-������>zE�������M����:�Z$
��~c��}�S�4>q��0N�����;��.q����ݪ5FP�} ��y��o>��L�Rv;�xAF�1ߧ�<K�PR:�5̛�S��]G>
`�Ő����A���� $���l.N6]:	�(p�Kd�Hc�Q>��/-�2w5���D��/�ؾ$ڵ��E+���D�b�Ɯ/C|�.[���t[酦��z�����x�!]���}��>�RF���.�&S��1ȗ�w���h��fϚ���"�<�s��'�ky��+���7�ֿ�i�m���>���#�)�d_k��&,��c�Ot=�g�w�U0��{�F�pI&�#����9/��6���z{��`4�vVŠ���t%�ES������4E3[���J���r~4�t�7g��O��,����⩝ޯ؎�M��~�v=����M����Ov����H�!���B$�o�}"���LɿhXJ���/��d@�,��{M���E,�jb|��R��<���Vm�G�·�%��[LC)p��LѨ���!QƲ�޲Y���8/�l�tA� �^��B�Lҵu~��m-.u�G��@s�x� -�y��̓�[����"�j��[јݓ�mR{��t�'�ѕ-��{�đ���lB�ö�n7���a����s<]�a�W�g��<���������h沸��=4�[r��m���=1�7qxRT���d1$��m���K�(�#o�Z1A��"\¶UZ�)e~�_B��Z?2��I��¢r��D���Xoj[��p��@G'�݊�#���4@��q�[1�E��Ki�Va2����;��E�Gxv��Od5	�څ��uu�����k�^uPG	>(]�}hS]��I�w�p	�2O��W�A-��ɳt��N@�b��v�����G�q�w�ݶ����J���=FlP���+�e�P�,�I"�F׆��0��;۪((5hIOQi��P��7�D��h�F�j�a��:��U�2O���}#�8��O��-e�v�/�\_0m�Ά�΍u9�
q]l�����R�݀Y�P�TN�S�~p�i�Wn���#���Qd��r��r�Vl����X�Bŉt����Q@(�����z6�Y
�Aj�����@���\;ɪ8�V����9S��[X�L��yv g����d�d/��>�k�ͦQhI�|��?Ϭ�=|u}���ݿ�~A�o�5�ݍs���ɭ�������rfd�*�;7��C�<$L�wk�܃�������207�Dq��.��V�K��/ו��Ѿ���O]��^����T�_�z�����*�Uvu�:����o�{Ҁma����gP{3�@V�Ͼ����+Ō�Ѱ^������Ď�Ì���V��}zK���r�r�{�AbR���%[�|U{0~�E��f$�č�8{OXcMMh�:� ���v=�?��&ݸ�f쀴����8S�Q��B/��k!��KF��Bf֚����ֺ�����*]5�c#���b�'a�X�&J�X-�7��Ƴ��{�}��ԟ�=~>�d),�=��1�H2����XM�`������~�s'�g���q��e��/}�~��7�{��o���' -DU��$9y׋�����?���o4��?PK   x��X`"�v�  ��  /   images/adcf2c83-f38d-4d07-a246-237caa0514e4.png��wP�]�6@T�D�ҋ �Jｷ���Q���7!@��H� �K��@�p���y�8ߜ��f�;��u�u]ko��4�	�  ���� �� �߿�����%�A�d� �)`q'˾ Nb��^��g,߳4�~�8:���1h�xnh�����X�F�>0(cI�4��@�X�&X��撔f3�n�K�`�I�~~�?2�����5m�Dr�L"�Ĉ�d�q��
�RO��R�j�
�/�����{\�[@mEE�Q3!�U:�oV�FC�###��/�x����Z�Z�%�2�qr�� ���#�W�a+++�ٿ�����! �n��/���� �T��V����9K�m��~���
�=[ߴ�����ݏ�@�l��h�8���d������� ���1� �Q���<qI�_�$`�qaw�Ϸw������8��45�����U�����O��� e�UWW;sn������4�8fVc,��7su�2���3��$��ŵF����۬_d����K��J��Ӏ����?�t&%��~_IKw'�9h�E|��v�ٺqrY߯��I3��2�+�l�x�`t�{�WgW�p8<��=�~�W��8��ܧe�3cz������fۏ*7<�W�̎���_����t��b�y���^�(��ab]h�wo33:���L�J�����������d�s�cK}��A��SOȲ5;����y���ƙ�xf�Hy�xn˪I��UJُa�X�<��HL{�����
��o�V&��0
s2*Y���b��犽C���R�܈�MaST�&��/��g���	j�ݢ��b�)J�Y�2ɹg/!c5�{�o�T<���)=a�=��z�f6��=�1"ؖ_���������U@	y%f�.>��H�c�W�˟�m�z"Ǆ�:�P>9\��9As�MRd.���k�N��H����Z�G�y��8�����ގ]̻ud 6��i�d�SU��l�G��`f��ȼ�LO�Ie��O�(b�^`>���̀/.}k;��%��7k�O����0����5����� �#��y��U���-�_nq��05�YK��<T*���6[�t6�!�8X��J6�Y����;<����l��6DS&�����@���Y~�Rܰ�%(��8�x���I�
�A�lcZI`��O�7Q)v�]�4~���錼�Y�TPY�Ek�n'OێvI�doD�_�I*�	�w� �XeL��,��l7�A
�PE�N ��-�}�m?�Ѱ>���31��tj�b�ӡ�~p�D�������MW��g:;��9�<�h��,��E(Xё~M�$�-�n�Pq�Nv���8F���԰(^		"w�T��I���_<�Y���e�>7k�՟ �h<Z�2�?c���AtH`b����B�e5��˻�s?�{bS�x*���37G���`�Zrg�qoM����)p?	��0�w���y$�!I���h5��]�IH�!Q >੐*��8L��s���� }����/"/W�;U������w�?�i�~�z�gQ�����\�:���OE��X�ﾏ*�~xT+�����]&]�^�Z��u�W��MG���=���у�8�Kܦ/w<�|�;��hP��_<�W~�Ҙ�5��\������ƪv��ϒվ|i����Y:q�D �Қ�daK&�h.��.Ϛ���ZP.^��1�u}�����kYa̋�y�,o�]%I�����C�|{�z�[��s�o��E���֠���xI>n��)�&ҭ��!Q	W+��D�V�}/��/�QY���������Ԧ���Rջ����y�.v��78 �IF?�[m�Q#�G�%[,��r�E���I�
��"�Ek���0�����:[�;�nb�~��2�123R�wǼ���g�bQf9�S³m���0�L��֎]H�󱥕?U�*�= 6[��7�-�H����O����o{,"dHb��승��f�qJ��.�2{�6s��K��x���i�4��~�%�*��ff5PJ�\���N@���L���(ͧ�0L��ܳ����s�g�������K�W�X�|�s�=5�]|o�(nݟ��1o���������������ڇ�=P*.��$�2�)n�<�O6a�$��έsW�a�L~^<|�q	���Y�ޤ�K�t&��a �w
�����R��9�\�e,R���h�������b���M+ToL�H鈠���t��I�5� �0Ǣ��R�G��g��xIV{Ȋ}*�7F�U�zv��S�Ƃ=X�����Q؆gk���%o��>x�)6�xP�m��0f�Z���.�u�x6��]9������`qw�d�����X���u���m�3i>rϠ�U�π3����g:b�<�p�d�,l��q�
<?](f�5pus12�oS����)�܃�c������s�#K�����7E�<:�j���ݣ���d�݆5��6H�י�=nRY�ʧH�r
��j��o������
+�By�dWJ��b"�3H������@�DA�	c�麒18�Rc[��Q��v�"��(ʋ_e&h�V��XY��o1�u_�[�z=���Mf���G�||�џ�����%��ixz��p�uA����]�����X�C��R�gg�%R7�ݛ�;�F�U�<���rf�s���yd6#��=�$���)���Vs���6�����bP^��˱�y�mI�g?�{j
�Qi�]&�6Id�2?_���X;��z.���u1f����)�̛��fAZ�RE��ěߏ���n۵Q�e�$�I���@���mn�K��֫w����Պ�����Ю�7"oN�i��w�!}��5(&(��N��
O�^t�V-��w�t�D�h�0����Cy��;�%Ò��v�>�b�K=��-z<�o�C��~��9LD�U�qjѢ��n�h��i�<�/��\�����v;Va����l��w�)̵d��x�&cN��� ]?��Z���������l���!~�[q���J����q�9�Iw������<a�����ؚ_���ޮ�(V��?��8�)h�S��'xx�����HJ:�#̞f��w,c1o�3#��c�Xה܍���48��w�{�Sh�v-���Qq,g�%;���(E�(}�$%}�t�y��5�)0ٶ��|b���/|��0J�p��m�噈������j�h�!,"��<zy,���QV�uēlb���t��W����?����d7Y&n�>�[1�in���NCo�S�ݭ��W����u�k�ol*y#��メ�8��հ�m 0�M�8���ه����q����Xf��}�F!&k4�W8�d���?�����r�C�p�1�ŕG�G�Ȏ��<m��}s�����'4l��o�{v�W�.4y�3�\�ϏK\�����j��xD��*��dqWb!һ����$v�C��ն���:���}�]��)a�������d�yI�}X~�#���@���{��PzY*E���"g���{�h��/g���R;�̛OG\��"��͚|ܱ�,�ey�%|�̞/���[Q>q������=�<11��1���=Mq.���	��j��Br�VG���^�k9�R���!h���c�ff�ާ���|�x����N"[��e�Q��Ϛ�ݏo��V���`���X`/��c�p4��������͍�֟tgۯ��ٟ��򏐚�����w�����$�8H_*�L�7]u�Y���)�l+���.�`��]ٛV0&�%pr��V�8���7}�Oԭ���4t���4��tmL��}�V�ͮ�{B>�P�ZDRr'N��K���,E`����а�R���6tv[S����_��Xɫ����O�̸ 5�w�.MS#^������q5+��D���
��6���T-�U�(�q�$�����yNh��܃�d��*�$�AjO��b9�@JuQ®���񅋾w�L6�Dp#_�n[}���� �T3Y<��v���ߤ��/�.'�E�J����'�l�n!1�J� x�"QY�v�솾"
�x�D������J`1j?��dɇ����4aE���Uq]〕� �����]q���A�bl`U":�~L�8�{߮$�0�]�(�6[&�"mi�p��M��},q�߃��s��y����/��t"���T<eA�a��/�e�������M�U�gV���2G���u����Xޒ@4���a��~�_4��+���%Sa�a�?_�'ŀ��e�Rb��w�*Z^�*��S(A9��^n����H��>��>�& I���n�*��/d&9�
µ�LZ���Q(��j�c
��ǀe:/�[�Lu,�^Z��k,T�����8��7J���v�LaPކ���X[x�7Xc�wn��^/�%��(gˠ%l�t�Da9M�^:[����~����;$i4{уن/����25:^���*�p�f]�Q����_��s�:�pd?�l3���rw�����8_bE���)p�C���t�nq�La������)��кPmU�y��C��N �ה��_�B��x_�=���8��%_�<�^���JCy�L��w�PR�U�?yT<�߱���&��;�Q�ۊ�%�������O�{xsBb�Ǫ%��9mk0N'P����a��M]+��Jp� ����ޢ�m�8�Ê�r���`Ip������ş��l��?][�%�{tA�����j��>���1�U�8�@���U>ρ���v���e؃&��1�.ͪ|r��U�:_�%�,#1cܕB�%vf �)�qs� �G�n�%�p����ͭ��?�������Aj*���N�T�1&�t���Z8� �=�VO�u��ϓ��)r�L(�sY�$��_ c�09m���y�[���7�;o�6W���䟓l�@�X:=��$(��� /����}TY ������,\�R�~��Ђ��dL��{�E����j��	����eKE�|D�t�'=%�/Eu㕻a���,���F���%iE�X���L ��. �b`�@uT�?�����6)��3�8� jo͗qh�'�@�4�.H�{�2��l3I�ݖ�J@l�'����������WC�j�\4끡�Ro�Fe�|�5ܺ�Qf��b�!p��g�z�p�h�djX����;
��)%���>Ss@-iS���1;�k9��-kx��rM
 �G�L�u�z/�i��Ŵ� R���L�a���AȮ�l�wmH�Wͮ�iiYy��z?�
K�DW�܌6rS;���u�\>҄�`�Q����Z�Q���M{νWW�ۤ�5��g������=Մ�ǾtSIbt�h�ߓo������Q���;��#_�Qm���,~��W��.�&׫|���n� @��
�3EU,l���������U�!������J:.L�؇}N�4���b_�o��$	�$4>7��0x����$Cc�;Z�h.��5��o���������E��h0���;i�f�$��gb�;�4���B��
Rn���y� 3�$h+�_�Z��65�O�ٹi�}�����(m��*&��{\.�Wy!D=xX�l���P���L�/vx3i�P��:-w����bg�kK��`xS]���|>�;�!�xA��V:&�66u2`�@���$�_�L?U�����Ow��*L������S��./$����'r#)�Tj������[��ފ)���ξ/�F�i���Dx��c��W�x�(n�ӧ��jĒ�)��o��� �k��=�h_"
9@�(�o����"Ƽ'}eQ�ib0��/�����oǎ���#A�����;�b�zy�a���[�^f��y��)�Vy�)��_�}ё��5-�I%�$T�z�����!�_�ZK	0T�M��dK�L�=b=x;Lv��x�{�*?�P��x�c�&:Ud}��[��$�|E\V]���)���ވ=���B?�3����J��䆚��Q�6r��'��9�P�m��+L�OH+��HHi��<Zʧ��12oM⹨ZH��b���Ȃ��S~O2������s��o�T.}����]s�)��l�Ajj��.^��{��?c��p�
<ۨ4��;z��Y��&�t��_n\��5�'�T(b�@hM�4�#3)n�oHV+^<y3tɯ����}��˖�X�3�=6��NU��,�!4�ۯ|�r�3@�ƈί�R]l�J�'�{]ʹ]�QK/�����#���al){&��
v�_�ɛ�Z)w:^.���f���2K��@	~a5e�����䨂���m'���x������	e{1�3��� �G�`m�3��6��$��O�8�y"6�^�[�Xn�3���21�	�>6ȡ�B2�t�˱	���R��׆��� ;�c~�愙Y��R%��ח��x�ېU��=��Z2>�B���p��`�O�6���y��m,ۖ���ܠQ�X �e�|�71(;Ȗ	h��GN-�E=��8@=P˧2 W�wDm�w��FK{mϫ�z� ���g��Ӵ��63oc���'���V�! y��5<�>�%���鳘y���i���{�W����=��x��u�O�^s�>ӻ�4Fږ�JQ��`���c�4^�^��X�t����H.�m\�k��ͷ�C9ى��õ\7��k��=�}�)shz��mF�KҼ֡`�p�:��=sI7��\qzJwh�����%��ܻ���Q�L�Ո�t"��&��"d�ʨH�64-�!י����#��f�d���Vkq��eE�2��@��Ԫo�kdll9U��uF)�� 1ʉq݊W'ei�ɳ���n�l52E}6��D���Jn�yE��_r3�e&S�^b4T�]���)G\�6��:��c��Tm��3�[��A���cG�8v�^pb���Q��95�����=t��� �ƇN���N��<C��'g�W8�^q<-&��B�����s�O��`��_���DN��%-��T�+��0B�ϡ��򛹦��Fm�����N'�-���Gf��W����e&";��ޚ�w����DҸ�H��g�9��x�C6#�~�ԑ���R6l+�O�?~|n� =D�.�*?[�n����AV�_��Τ>�6�3� ��	?�_�Q�!�� ���DJ߳�Β�=4|Uh4KB�๥�ΞQVT�]1+$��|�J�N��	ߟ-R��L�}��p
�k�=��]\��<�8S��I�[V���в�W�a*ך���KY�2?�E�!�7婝\k&�S&�qD���/���Uۈ�\����D�G���kb�$�y/�[����F��������ń�^��7���8}���K\�%��2��6]�����sƞ6Ub&g>�مB��T�9kz�m�Z��zE��T�e�k�������^�V/�5�0r���a[�)�"���A �q;��
��[:��(��U�E1I�D�M
��	bS|5oٻ���A^��66�}�"Vգa6��Ya6�A�Q�hF���8+��1Я�Z*3d?�f(�ck�6"�cύd���I(��{���!E�7��2��%9���J��
t(�G��A��M��`����ŷ`f[l�O0Ì�#f�sq^���ggPܩ��+���fy�+!�qm��`�ا�2�DT	j=Z?\�ь �����Wz���/bB����#{wN\cU��l�`�D���[_&g�C�a�y�U��,0M�':8(�q�j0+�ڰT�6N�_o�a ��� ����*Eh��j��"?��A)�-S~���8^���>-Q�R��@6���H]� _d���
�� ���i���v�^�u�G8	���^��7��(^i�0�����U�j�.q[�*6�6X��.��Ϣ��N��Q�i]�ϟm�F"~j�0mK�FĶ9��B$��Ը9b������7[��'s�� �Hۻ�W�l���E���#_�4Ab.����}}���l����3�)'����g�)�\�e�|�8=��e�����	/kꨪq}�>���y���7n�1��(X7�I�0,:�(�����55 �M�?�e���Z���/Y������j}�+�نyt�쎷�������	��UYW>)^�[��&����g���t�F���{���Wι�Or�Y��Lä�xP:�%�g@TM�u�:ƉXX����B��׽#��`c���	5��u�(1"�q�
�y��E�i��0���u�d7R=�^~��[&����`�Ԣ3���J�蓏���j�ڴT�"�}Ϊ����]�W��*��O���3�Q���������F⅕��/u/H��U.�3U������ʡ�Q2�L��˓�U��+:����2���m��t��#������})����� 9�����霜/�T�`D
�H׿W��\'�Ф�՚���$J�JI�eh'�21;[en7��u�p�&£�l��p�\B� �҃�/�*����.�3����ߴ��>v���q� t`�w�j\���w��u*	Wn��U�`��O
�硨�W��RӚ4��ܲ9\Eή��恗��A�����-���m����T������E����Z"%JES�o�-&N[�z�M��#f_�.KJ+uD&7|�����ҕΎ��M͏']dd�`,��W��k�n��*����t���K������Xx�l�1.Vv�+'�x rwE�޶��|��=�Ww�[l8�e��G���nWB�� �9��h�����b#�R���:Bo�I���葤������Y9|���r�˱&G�
O����!ׁM�a�͸I���T#�F�1��f8�0���m�T�Ha^~�?�SXb
A_�4G �[L��̟=[��jF=���<\��i�Bt�����uJ��:��>�y�Zn����0�����5xf�X��vj��(5y�If�Vf3(���}g`�@.F6���MZe�
�\#���)���u����;իņ<̫���q�I���Բ\��77�@I�y��L��c���ȓr	�wC/��D�bc�'��"ΠεI�{�Q�c��{��������DHG��W�S2�IހȰ"�q�� ����̕���:8�>0(ME�!5��/�R�	P��,@�oP%�rrU[n$�� :�=���Dz�3U�
��#-�|���*�s��=���8�Eڔv������n�����i^fP���A�q�v��F)����ގI\k��F�c�������e��8�?;OM$-�[(&&sY�{7��6����� ������R5B=ʃ������bAϵe�qk��ZW���ҹ��-�t��2%�(�� *|�Z��s桾	�"�X35N���F����9���x�v.v!���L�sH5�]��N�w�`�J��4�� h��]i�G�?��v]J�*Q�5B��b��Ȯέi�
rƷ��ۙ�-����n�(C�!��o����b�K�`՚��z��i���z	���>>b��A��7a�:c裬�O0����8ս����P�w=��!.X���'||�B��8ڧ5�9 *.�^���k�&�O@�({`�ť����� &~%������� ���*���'���]VI!���� 6_<FGu�\�dJU�y����m����9���k2��v���B��ws�؃b��'��\���+�����f�4L!#�6��O!�ݡ5(��7=S&H�}��B�^��}MG�#lx��WԒ�[�2��
U��>�,���j�=�m9���J��
��~�qsv��)ZZ�'P��=VfC��t<��S���߫!�O��f����IRM�.%͐���
�{>l��7t|QPk���Һ�,2��pޟ��XZ���SQ1�,j51���p�X)rJ_�<uO�g��Px��]JD�+�x�Km�+c�8�l��^�:���V���-8��d�5���Lf(Q,/�L:ag��q$U֐��t2�5%���JȺ@���W��b=�h��Q&�y�_�H��>u����E����t��)ޭ�)sA��1S�B��>��`)]���Zߴ!�`��%�)q�s���N��]��m1�LK��4�O��1�<L���?�7�j�snu�eu�= }�9fS��̓#E�EWg��s�$sv1�=�L�@W��S;3��c�p J)�t��s�a��>9~�8�%��wD}��^"SJ�g*?���2Rπ�j鹟F��aذ̋��:?��0]����z�'��֪
��cx��s�9 i$��f��k)��ۖۡ�=�	��k�����E�Q�vZt����b�R�{7쭕�@�s�����7���mC;݊�*�A���R�RuRE��j��e/�l}�LE�];�I���!�uN���Ӗ����4�)+i�R��ߕ�����_�uwO]�cz�Lߘ$^�Ǭ��MHB��ܧU�!;�Xw���<��;Y-�;ޠ(Ũ����������8��?�	_	�$��Q�.4�l&�LnǢ�C�Tdy+�-?c�s��g�%q<�p�CL\�~�#�Z��� `�f���~>SZf���24�&��#Hq%&ב4ԩ�1<{�}L鹽Ŷ���q@ͅޭ��*h�ɭ��ٸYA��J�o:>!��y�!u�>�R���E���GZz�XȮ���Ϗ8e>��lj��\�����G�)�~y1Q�w鋆h4��2]F5Z��Y��H?�G��������7��,GJ�l6���窜��Q���{O�,~�O���U�Su�/W1��C���=)���m�]#�J?Q>8�����
~��	5y��?S����(�nO��Z��.�-`سp����/�'V���2Mv��r<6G�����8M�U,���h0�6�K4P%���N62#���O��z,^�r���+�Ě�ۮ�c?��e%oH2^�-`�T��\�T[��k�`����Ҟq�-.��Ի��G/M�y5L�k��Ǫ�E��n/�^ݭt2�J3�o�qE��v:�O8�)���u�=��Q޳��yY���9�� _S�;5/#��E�l9V
: ��
A^4M\��8e�'@��&:����&�F8?]�OA����@J�����j�e�m��ҹ�]��k'=qC����+n�F��k�ѩ���
��8'����K7RL:��^�s��ܹ�� ���DC����!���^�<rq]iP۵���U&
q�:�j<[��8�b}m�Z
_����u8$K1��
#�@��\%[h5�t���)|�uW��x�|��2�Uɟ�1����㳄c�a���'�ٞ�f�?�p�4zG��SF��Y��7�Y�s����x���'� !� d\��萺�{b�µe�k&�NklpU��΋/�8'�7�=��|ܶ��&QL��z ��$�L�'�l:�U�0�uh��].6%p��3^�b������h8��Q�,�����i�ļ/��,������{�?w�<Zy@O�r��zNtmWw��/5��B�+����d�*e.�$=?#_P�mKM��E[�_��Fj]H�5�A�"*�7�y����*��7�ʶa�Z��d��lm����;\�a^�sT�3W��܄��d��Yf�^��|^[O#M�Πt*�Hk<>�s�^�q�y��*�*�Xڙ��$y�}�䋧z���Y@�!	l���*�v��Eʤ��c2ɔ��?�-��mE�c/�Frw��Ѭ���s|/����꫏7�����G`�=��oQ*[aF~�f������۳5%#��:.���x�Z��s�%��o��w�MYP%��q�6��|��	|8i���]Zw1�{���͂S$QTvN�ǍB��9~�Ic�c�� �/�R��v�J�������䲛�)㎋@͵��(we����'KP��6J��z[�!�a޼6����B%����l�U�Qp|�7�� �����i`렫"h��J��,��G��W��/u(�Q��2�B*��A�ނq�Y\S�4�^�,�̈�6�f�-Cg�[V&����`�/��,D��#�\�|�UY���a=�|�!���Q�-Ǜ��3y��z�I��F�@� �a:ץ��{~s3{�ؓ,�����;�2�l�'���n�<6h˯=���A�܊��t��ت-�Z�V����W!^���J++�_���G�}<@9p����o�)��R����$$hP�R����U����;y9&WK�.]ݱλ�ʈ�Y��ݧXc���f}��D	lRxF>m�2�(���:]����VJNƄX��	���T����k��y��_�qO�wx���f�tN�
��>���i2D?΢��x��Qho���g�p�/۱�&�B�	���x�u)���t�����ʘz=�(j(0��:�-�O���[�Ժ��Y<��s�>7<��!��U]Tw+��)#�*u6���(�E��P	^�tHU�hłW�A����끝�=3>U�ֈ���'gW��>����W�bz�m7�6���g/��c��\hX����B���-�����Ë]Wʶ�l����Y�ϜqWV���מ.O�mD��_̕��w(��?z�y]��9�T�Z<������CQ3dCAYwߘ�t��EY�vrJפ�ȠAl+���c�zA��ǰ��9������$�1�|�M��1NR�U�W:>��뇡9ZGW��3�������3��p�0���3��l��X��`B�ΐ�<m�l�~�n�����L�f�A��|޽1��l>�;r���叩?�*i�2%�Ī4�O\\���Hm"
*x$��G����.�⥚�~���1T���^�\߲D��φ��N��0�r�r�8����N�CFg����Ēb���𘎻v�N��@}�e��6�w���!�5��������'i��\�IfՅ��yW���0�1%az����L�IQ�gW63K���8��L ַbR9�z6^g�d�M�%����	�җ�7�n;������D��o�Oq����_s�uQr����5;�<}e0ٹ��q(QE����Žx�}��e.R�[�Е��e0'u�PϏAL��<�S�f�X�{���ǈ�Wn����<���0���=�=������ΰc$��ڌ��hp��_���D����n������)�=�"�=�}^1U�!I�*�����M�?�܌ޱV�J����D���C���v��ą�/:�CT�\@�FI	�L����Onٗ>��WYV@<��H)Oգ��u�����a�_����ߢ�Cz��k/n%�w���vF;W�x�>L�Ǽ��F���d�.�҇t?=�(�A�ۀ���y�J�)�r&��u�v濺Ty�r�.C�_�Ɣw�z��#/���+���ɨ́��Z��bm�\��a�Oy^�t�4ѭ�~����I����^R��V~������;,�ދd8�YX;�����w���W+��=e��̕$���[�O���Im-x���~d�*0��ܽ8]0qք��2�:aE�4A&��N�fE��8�r��\S��K�m�8�h,�[Ivt=y�6�~��-�p��p��4�S�Ь]np��3w���
����!�R�9��6��ΰ�ccӚ��(Ɉt���dTL�@_�=^�����;֔�-�V�}t������U�����m,^=&_X��}<2l��SQ�L���C�aQSi����z���2�A��jg��{|�EmQ��8�@�Y���L�'>	��f�@6$򏛲6��a'A�HvSh9?_�fj-(�8u;Wg�;ާS�d��I�(�_����Y��}4f㌋��k��I������,���s�:���v��>F��X�	�(z.kL&2h��#���.7֬�RRb�7z]��E0�.�����Ki({f���ZCZo5�JD��7��-�р����?;׈�wY�>T��0.�Ќ5JV�9S��H�Іjt�`S&a������X�� ��ʡ�-ezB�����%����TK��������3Un���]�P��-�レ�n�n'rs�"�Tލ(p�tKJ�`u5&OV9g����a�kV =�Y�c/j�쌹U:�'T���x�ǌ�J��;��⨱�=�����tm��Z�:&F�N��m��&����4� ������)�$�N�Ȗ�^�����MC/�ɾ�S9���Ŕ�e��s���Ip��@�j�|��gV*�z�清�0���p5��p}�C�y�­�*�/$��F�6�����W0�er�.(`1d6�ӘO����?�Np�3����z��?�5�;]L�)���{9��/Ep�P���e�5��V	��I�ÛkEY�����j/��2U�#���9μ���4?�9�O�����Mj�j������*>C.J�(nz�h��$d*�ߢ����"W�u�)3�J3�ʏZ*��J<��E�^!��Tx���@uܘ¬d���L2q�����!xL{���`�.Z0\��*~�0�Т�#h1a��������X�du��LY$�T₉�a���{�X�(l���Q=��p��R�0 �,���4��E�;�]N�zY"��@- �q��:"�@i�m!��z��]�׽ƣU�N��/:��s�v�ʴ�|5�J��6{��]��cPuS���dr�;��;B�Ta����~��J��ؠD璮��,��@����O�ѕ�E�\��$�p���ʜ.���+�24^}��m�n�\�!��OIV	�����huȴȫ�M>��,��ܨ�Z.���SH4��d�ݹ�q<�I��F�R�7�����Y�eԵ���a;�\J�
��S��2�=��0���G�֭VI`1Vʻ���}��p���,� ��-�Z�yZ�0k/��>̥�m��m;@�3I�x@A��+�H��zx�������n��;�([K��gp�4A�o��E�E����i��L�"�7�9h����_曇Qw(�
��<;)1����
�(.	n �eso~���м����B��UKQ%�a���?NIZ0 ��c
�L<�������E�f� ����v2��P����o���|1�u#�����2V|(��ց�������oL'�K��Y<����A�u7�(����4�aE�I��bL�ې��j�|��7:�3������|�d���I���f~�~�?�媤��޵ڎ
���q�i�~>��Ý�Ÿ!����=8���
RK���+�yx2X&&��∗��G!z�$��c�@�o'�˝6�)�1J>��Q�!Zz��&��e��)��ԅq,�ߌ�<��3C��x���QTߙx��G�k\
�fFsh��b��mvi�$��Zzw�V����젒"[�Fz����;�8���RQfU�2�$E1�b�>�2C'��k�,�i;�=E�ZC|t��g�o�����e\��'���`�rۑr�3M����r��s�eϦ ���A��w�$� �$|Z�n{�RZ�c�+�5&����g�Z3�K`|{bʄ7_�g沢S}�)}��θ76U�ı�84���sn��U�����0�����H�@�f�-����e�۟��!/��qf�P8�W'�a˕��G�7;&�==���4S./���o�A�!����j�ɴ{��Ye���p�:���ca�J{#' TÎ���N�(��IY�s���I�S���%��[@�1��֐g���2VP~�eL�r.��4��%�F���X0����(���4/y4a;O�V1
"�V��z^W� �a����4��ӅHWwp�vm�2#����4���4������p/��%�Jz�>��5B��Fl*7��=��pX�@�fƇ�І�W`#�vY���5��^<-����휂x�/�/Ϯ�wR�ޟ#ͳ�A���j,6U%��iuܾ�O�ˮi������mX�D�x��i
e�u����nՌ���h{c���@U����Qzz�-�Qa�N��4ľ�4.̆-����=��&l�L��s�Ft|�b���r���Y J�A-qva�$^�.)?pu;!�V:�M�V{8��������ˤ��J-NQm�-�pMM�J50p�2pKq�3��l��{O����>��jDh[@�MXƻw���kc~
�v+^��l݉fbc�~V�>���֞���{��A���!���b<�J%99��}������.};�ߖ���	�έS�/8IwhW���r.|�%�y�z��@���el�L��7�o���r�W�|��6��u/h)_|yQg5�ܹߴ"x6�#��7��L����z��b����L���ښr�Cp~��?W!����ܽl�1M��������(�)�ZV��1$�2W9pj��g$�u���۝r&i�􀡡�d˂<f��*wwg2��^҂n�)���-	�O9�э�7H��H|��x;��L�*w��4���aX���h�C�/��뉷���1>����[�3P���}L㖒c���6B*4��K���o��\<b�U9��~�u�X	;�Uƺw��Ǹ�J���%p��?	\�5d��U���1�RF�t����l���r

���U��"
v�������M���>����`SI��x3h�8�(�X�h�P��tBE�{��������^T0�pO�NEa���lƋ�y����l'�����1 �k�y�g[Rx���o��Bfhk�_��P^��0�7��ͬ{�*�KSE���I�W�!��=̏u���]���?6�
�J��������-'�J$������˽�o��'>�k�����
��5��(N����+r9j��͗����x��nr��|�r)��/�~�KxE犍�a�૩���n����{�x�ABI�.��.����i���a 鎡�;f�����|Ϋ�߹�^q_��Z��x��N��o��T�,`?{��ҝ�ǻ�	��osI,��yH1��_���nZ�i�9��=(����֐�O(�B��*��'��Z�ZJ����e��m�r���ظѪP����B����DuZCSo<k
����"��r̦�W�A��r��k�]5m$�����h��҈U�q���_6)��EE�s|1��멖ߍuˁL���;N�PƧL |����;�-�nGN��h��bԇ׏��0�m>�ڟ���Ηh������	�����w9���D1�?v���̇%g�|����Zi� �Y�<��S�\��##��q�N1C�
'���D��[�hdb"�KO���U�
?[֟�4J��2/��)�/���"�^�,g}�������!���h�XZD�|����ݻ�c}���!^� :�=tG��akW#�&�K�=r�͇z�gT�2<�
N)2RG���O�ĘL�Y���8`�	��X𒖓sa�zpԳ�].��:��}��*�����+��X�K������B��c�Hx�3b{Mz�)+Y���ʘ�D�G��6!]R�X!��,dz��4���O�ە�`�ۿ}[�]:I}��
rL/.�a�075���S�\�3�R�Z��ڸ��>O��}���-�p�^kk���ͬ��['7Bx�ァAoe�ރ򿇤��v�unR��RaA�=�Pz_hԒ	|Ժ������J�)7�0�MN*v2��J �0�XY!{M�&c]�,����(�6M�(�^S�7Q����Y�>PX=nhD#�Sp�J0tdf6�P�8]�D3џ��~v�i�ٰ*�U�Zԯ��C�2�|k�򲊆����*��ǐW��T�����B#�Z�f|_��#J�I4H����/�^��$�D飱���R�8
?�����S�̝�����<�K��J~��~�'�h3'<�����I�U��?����+���E.�2��x�U��sqߜE=m�-�w���9�Ռ)�`u3>G��1Եw7���Ҟr��wg>��s��M���]T�D�h�-yZʙ�.3�t���(��t�R�����L��AdZ�����7�H���KJ@��`
��~�I���:֑K����Ag�`Q�) �or�KF�������?Z#R���'�M|y��сB���=2�>��N�pV�	����=�'r��Ģ����3�H��Y�}lm"���.�W�=�����ʻ8�v�N�'�r�x�]����� 
0_Y���8)cb_:�	�Q�<AB~3k�&q�yT&"�w��k�Ix��n���Nr��.�����MBK̕`�Bᑼ@��>�k��4^�� N7d�]��� 3?��Ce��(�����>���.`���E9b�s��w�pu����u�����R��^��mC�OsΣU	�#֑s��,Ց�[Ԓ� k��{��E�xD�Z����ƞӽ2m���v��[��m�PK6��&�� �P>����q���~>���8��O�_3'��]:��M,J	Z0H��#�dy���S�#��<���Qec�U�u���pӂP%ˋ�E�����*�7�[Q�j�k�p��f|�	�@���-O�B�g�҆��擄E���H)�t���g��(L.�"�RKE�y^�s��+ {w���=�s�?u��M��[UVc*\��.���գ�	(1�=�x���˨kGS>��ʹ�Ӣ`�r8�&���	c! 	�C$5"zc�ol��i��s��{g�8��3.3'3���0�����
 �������n=f��&�8]2_����CήC�AȚK����г,�Z9��D�f��	=��Hnܴ�	GVz{�8eoO��fx�y��h�#*��)�n[���f�!�[1,�8�?BVѭٵ�:�}AO�l������\�@�x���sR#G��ce��3���$M�9UC]T�u���=$eC���g�[�h�Ըb��Z�}H`�Rl�W�cV�<�:��~�7�&�J�fO(*Q��>*f��r��L��� +�!��s���p�do��-�MR��	u��tEfD�H��~��껌o��sw}��=�/m�6�
�n<�m �T׊�^�,����Z�	-!�2�_u��\�����R�?T@���C�}���(.7�<n���@�O���P���2��g��J�*��2ϰ��;���1�t?X��N�:S�]p�,����P�Z���h�n��y�U�������1����k��n�Y������I<Gh���u�5�U�C���H�Hw�`��%�
k��E1t�c���#Ts
��4��L��ǏCqx������'�s��~���١ӵXY����<,4�y�q�ۊ�C5�÷+����n�q�6	�[B믃��+�<����[������E��]�v}�M8������\����y+e���k�3;�f�b51ݙ�f�p'� Y�#7���0ņ˃ˍ9ֹ���W���PT�M��OV���l|t1C�OWH	�,fg��^��t����g�{�|
Ҕ.�q{��ӺIM��j<Im�^�8��i?��JhTVj狠E� չ���U�����Z�+�����u��]}�x�\"ɇ[{� �|���9�������Lr{AD�e�����m��Ye�1�40v�g��`�<��k��a�Mq_�A�(���"��S���qS_�ca�w�t��q��||~Tl R�mNcR��]>�9�UWL��zǖ_��v��pc
��)�On-�O:��Ճ$�ye�>+���sK�Y}�xf|�m��H�ܒ1dG^�R���vk�8����JgW��{��L�ثA���]n��r�^�؆iL����'��A(�d؆M�?�;hN��]CTʌ��J~G��,c�Π#@D�%_kǅx����X���n^���bV]z�6ɤ4�������Y��@��]��ScK�R��]jh{����a��OW`�ZN�)	��է�O���eI��~1���wq�a������#P�{Nn�HaVq���/g2H��g.]I)�#��ѶB�W�&t�L�Wљ5�v2�t'�)�ڧ��h~<�p�X�z.Ӷ����s6jJ �g�#��$��Ts�zѕ��r-S��#�P�ٔ!����e0AEBY@���t�e�8I����R4�:_1�[�? �*~���~��dF�/v��9t4�:Ρtf���eX�e?wqُw��n���nįW*�0��t��1�4���L��O]�l��鬾g�܉T��XD��4{����afƤ$�h�ە�C��	dy�8��=؈Yv��ܯ.�����MO�K�Y-.Ά���G?�ls��M֐��(:<�M�vmM�8�H�n���		Q�7�r�d���^���ѕ��S�|ʤ�<y+��Y���������V�6�7�`���AX+�R�J O� ���+Me�`)?�k(>5��9b$�펄�ք_|��,���K>��|_�	v��Ϊ\�/͋'*Cm� ��D��ޢ���L�	<}��(><=�/��˩�==�Z�|��& �0F�ޣ��_-����� @5�*��J�-�pw�f������y�������ֳ��!	�c�##�k�&��"�Ϸ�n
aOw9�*��o1����fA�GF6�V��_�����9:���sM���9ا�.�	H�@�s�y���s��r�^�A��,�is�t�/$�QK��e`^�Y�\��;��U7����[��{2��y���RV2�4�W��}T���u-b.z�����T_�F����<bގ.A�Iݰ� Ԅ���L�����O/��O4��d~x��'�X�� ����u��!��No���S�t����án�eB��Zw�O�ZX�Q���9�+u�5�]���lbϫ�t�є!�I�d��.�����W�W�iJ�m�_�W� �zk�s���Zw<����ޣ�����r��RJT�mS���x�����KWi��C�����7x������W�Lz䂏�!�o��ˍ ����Z����L��I�T���zj��%��e j��8�'�l �2�,���dyhrIu��$]�K��_:""��*�3������s$ v����<j��ޡLOl��:�����d�����Н0[���,f��6(��'�Aw��idWh���R}�߯�O{���
O�F��E�APA�'���(�T
�?}�� K�T���W��K�zuG��6[�K�Vѐ�,����p�K5F�Q���)~��!�������5�s���|*�G�+yB����}4�In�W��H#�t�H��f�P��T����(��t���N��ʔ����hA;H#�� Uw'�I;#�00�����D�
cy�j����9��-y��8,��Ȟz1g��1�DL�j��RjIDziī����D������F�w�\Q;�+�j8�����4���_�p�����XL/ܛ���ԓG�����w��d����U�I��u��C`�ǈO�?�%3�acI�l�D��r�����%����o=K8i�q�?��2�z@�/'o)E˰�@-#��LC�OE�aR��2�n�Y��5�a�T�?Ci'y8�Q���Y��kn��㧔���V55k�N���DcM�\d�[�w~�$�0v:�dԾ��&cʑ��A��WMBT��@����	\�P���
��_�y>i5���'ջ�92S�V�}TU��>wC�б������u�񀄖 �.��-U�3Sm-$���� xe&�Nna^�DI,�����8���-#[b��_�܄�6vTmd{���M���UP�ѺU����¯n�w���6\q&QE����JaǤr��(�H4�*!F$ub��AsY(k%}<ÿ�zC�o�<�� �ɱ���K4�B�������,{J���`ݔ����Qy�Kފ���%�\�P����1����MZ"��CV�;! ����J,��3;�qѾ�>s�r�
-���L�\�p��զ�.�tF�T0N��1�p���Tx} $F�������-9��27�s�չ�Tr��܌�v��/�4���H*.����?Z]�65��P�J.�H�u�"�X��̪���Uw�`�
�~�Η����b���8M�-�����*[��"��=�����_^Ul��?ZaD�Z���sܶ����F����O��7�_a�;��r|ˊf[�� :�X�Q�E�Hc%𽫨�GV��9z?�`q'�;_n�'�iQ���m�����u���PC��BT�-���Z�k O`q��A�{ിBkQ�ͼ�|�
(�I�a��u��&��p���?hJ�m��1)�	)Ű����w��iO�V�ȁΪ`K�G����0�CH���T��	�;��Cp�l[R��iL��T�N�A����߄S������?�τ��t��E,\���h���4�ﶇ�B�̇�K=Ƽq`3�8bl�w7rS0�^�6?&�B}Q.�)�J�7%٬@��ie?�����O�`@c�OHo-L���##��2��z� ��P�(����
�jסcj}P,��@�*�j\$��<�).!_��ɇ��UWJ�(E ���_�Y�Z$�8'�4���ܷ�>J�÷1��'��+֕�F5����F���)�>�P&l��l|�xz��Y3��H���*뾾�p��ܴ��3rmVv�@J�4�Bqfl�Nr��].a;�p�/d9ػ����RM��ՍG�)i��q��1-� �t�zq�-�<�5���O�ة��x7��Ȗ���$��DA(�y'��2�p������O]Q���i��,�>#%�;q��Ǳ�Q?�`(�(}ɂ��3�g�fBxp���!ߊ8d#^6]��ޱ뙞+�b�>�3���W~�"�a�蘁VCY?{���eZ��ږ:����H1f�9���!����[ЎoZh��L�_�*v%3�y&Ұ�2��a�;T]�.6�=X�&�y�͐�����8V��3�w��ECI��i �����%��غݲ �*vU\��	D�A����},��]ZRz��o�o]�1���m*�h��� ]�&5�§�b�3/C!��Jx�Է��/GP�6�� i��%��kw�{�e�fA(��d����*�v��0�&��@�����
d�W����p S�֯��6zZ�]������UG3�5�߮
 ��O �@���J׋P1;���&��z
]Sb��79c��H�R@3�m��JS4��M�a�4� ^4^�?�_�^/�~�z�%�]4+�T��SU��2����j�Ф��=�h�A�Yo��p�<�.�o��r���+�Z�j�����w�ƹ��j}��腖&�؎���D�r��vd���`�M�l�-JI������{��n)����x��w�pU�i�m��f���)n�uև��j����>�<�4}�Z%���~8XS24�~g	v����Q��&����=h�ק(�E��)��{[��a��3P�w���RS�T0���;�/��5q�qp�&�8� �A��_Y�0H�J�z�A�9��=f�o���q\�_���i��3����IÁBԡ�����s�C�-����"JO�1�u�y�Wo�Z��V��(8*լ��W!y��oS�'D&޳�CO��(ut�g�I��t���K���vs�Q���<а�\�{|L7ַ�[��;-���	N����&[ps	Tק�O�y��al�e��W�
��>��oI�r`�漟��Gv�KGC����8�i��X���I@�R�4����
�n�3B�o`��]H6Z�1R��L�Vt����]�]�)E���� *�3�n���� �Ҕ��r�c���/7����ۻ'8�C\���[ܔ����Ze�xX��n}���Ҿ�|�=D��Z�_`d�@��3��.�B�%�S�7�rN��Tj)G��`$�{�j�?R�4*Τ��9K�~���5ﶹ�#׏'��ġߓ�mճsC�;Ӣ4c6˄��0��'iS��@�ǮwH��I�T���5�òs���vzE��[�h�P�h���K=����w��o��f�~j�T�2�?��PH�'C$�����=\�.A�l�a5F�E+ٺ��E�u�b�*���_w̲�R*�He��0���*��Hê/�[>��6頃
æ��tPM1O���S�USZ�i��
ҎS�����>`�..�w|��F�#�Z��Ls�/�6ݶwX5�+lJ�U���[�a02eB5�SC��t+/�h.�=��w��е:�f�w�)=�k�s� �����<���INa���R�e�-��^�Uu�O�[O�]ۦ�[9V�G���VK�O�UOޖKά�u��~X��w?*?u?Z�ֳ�b*��	����t=�#E�܁�\Cشb�
$e%���Y�D���[�rW޶]��A
�;�z�j��Μ©�دre;�BԔW�B�����]��m�D ��c����(Gt�"@��J��^Zg`|QN���CPz��I"Ir�*׷�-��'�t�>c��#0$��sl�դ���ܱ���\�}�~]�
��}=B����	I�@�\�Tf���임��O8�4�Ꟙ��[R��~+����2͑pI0L>�j�#�mY!j�b�ib�Zd���F~*V_�o�����c�:���/�^R&-Q�|be$D�n��@�gT2׮ ��B�pv��}*�~iu���6|�9�:�߼[Y�������&+�eɸgx�4�~�d�}ߙ[�1��{���a汩F;c�Ŏ�K�B1�9���U�c�K�b(�&d�������!kH\��7U^�n~vd	�u�����>du�����V�k\r�Ī������;X�����)�|�:�ۭ6�?Y��������#�l+��k^k��՛8X�����q�q=��
.І�e�T���JF��D<g$|����<������w��luE�6���T���.�Y�AR><Z`�IF&&Z�k���\OV��x|V���w������ݠ���)Dk��R�qm[����ש6���Y*�m>Xl�D���Q)�vd@<A�/�-;2Xk�J95/���X�l���R�
"���V-�a~M�ʢզ��:\���]}ݕx�3�J�3O��O���;,g���ePV�JTv�`ee��
���G0���b�}T �|ah���#M8pR��1(��vk�0�L��ĝ�LD�����}���(=�)G��g��HQ�����ޘR����� B��j�GQ�
ܮl%��~��#0���v��4�fƥ�D��Vd
�мI�t����3�ɠ^�����@|�HdS�
��)�oCs���]�3��ψ��e�7�"D�r��G��޹3v�a��D��c��/lBrd��~*wDo3�c=6z=d��u ��J ��A)6~?����j�o|x?�P��M�W6.7�Ϧ�@��NBRC�%���h�;5&&Fi��IK�ŉ���H#�܈tN�g�
M%����$&���F��Z�*�*���Ua��J���oc}���,@F�i�ra��D=����-�}=-��NXEDE�\d�W��(J�hq���X��"H�O��r|���Z�@��7%t��Q��}W�Sؼ?�C�-�C����
�T7��L`�3�~8�+d�Ȱqm:+9�-�yQv,���{o눶>Ǟ����E��q ^��1f�AY�5��`'ǧ���)������J[��jBS<X�d����ұ�>����Unu�M����(UΡ-�v���g�>aR(jΪf��ʉ��C�M|��8em�^p�h�o�/��Gg�J���[�ȴ�N��,Z��J޴fjyj��:����<��e�n���Țq�pdz3��c�8���ZgW$&��ȏ�9��Q�e��]"��B�^�M�|c{�Bmq%�Xc����W�~��n�d���kT�π�]�7ᩕW���/����Y,�1'`��nۚJۅ���7�A��?'��yI=<���(G�|	�06���a�8y\�r?�U����{��2�6�뒟�Ev�,��EɮO�S&`��[8��a�F��E)����C=t틵��ơzƗ�zXDkk��#�˟v�W+E9��=F�LOA�-?�:m���!���_�O��hE��f�z�aLU�T8����RT�0l�sq���r��JQG׫,6�[�8����I�3J~4JE6�nJ��E{I����^����[4������.��K�^�S�D /J-�1Y���O�-Ϩ����|_��Q���Kb���g�&��Y��$JUh\�C.4@!����k�}���Tj���������F?A��N��PK�Ŧt!�)�щ��.`�$X���ߎ�pמ�q�LQs��ȯ�x1i��$�=�����w/�c��M�j�H�Ve%	˸3Y��ݟ��>�3�u8hQ�W���x/��-Xw���o��}�T$[�_^7~�b�v?��/<8V2#�j�R����f�u�=�W��c�dsFL�u�"p�~z�:4�$��g*�}|��c�Y�h�'�yF�mtKcхA��ɷo�S�nZ`t�)��o�re��y�|O�B-)�Ψ��̚�3�d��ߌ�C��~������e�%�YB�*�m�HXF�����}D�(y���S�P�+|*;V
����Y!@�CXϢ��퐯�O8�!�9��o-����wUGjԹB��[u]d�!�m�Y�_�^e��s�^���diX�d4;15/�h���ww~�Q��BO��S)g�}{ �&�|�|��o��h�am�J��s�>6��1'��G;$~��N��i��L��<Y+��=و�k��J'�f�Wf�7OCjKl��I{�������� �/)�d6��F\�v���lg}��ꇕTp�t�8qS�hZ�������~���ދ���K�i=���F�O�����*�E�����c�����z,�U�"�Z�4.�oe����9/�h}��-J-0���oy���Ĉ��eBE\D�kR�	��v�\�;�&¾���<z����q��pz�����e������Ԥ�B8��d���'�0K��(Ymg�X��ͰkO�X���ί�雍�'+$l�)���*�K��z��dMym1*�t;�{�O���!u�9�ƿo�V4�6]�4�9P��hM�'	���IO@IV���-���k!���ˑ%����/wO���n9E�@��Ց�M�9���FG���.�+�p��J%�ט6��z0j��}je���r��(�OJ0B]�ǸYy�3"��r�D^���e�/V�6v�)��P�K���j��޹]=޷���'d�]��ʎ�~G�M������Z��Ϻ��#X��I��hO���^�c������k�`wW3��`
������B{; ���nd�����7Kٿ�6�[l�F��$ԑ�񺖿r~N*@9u\+����S�[�lV��8����� ��oyvp"�yI>���~�ɫ��{i��\�9���Cȉ��n�0W�R��:�Д�_���,�Ë����ޟAQ;�EY0��2���7?@�a��岐D�t�>����%az���މt��nA?L=�g�i^� �RLevפnQ�<�J�ѝ�N�T�����(�{�ͅ�Iع��E���(i�ע�fx]���D���X���]�z��8�u� .7{������<�Ұ7������,�'�h�Q��G�~��^<��!��&�Qn�
pca��.���d;5�H���I�b _(��"	I��y@��m��Ooݘ٭
br�ݚ�<��[�%�Z�yJ������}#��`c&�.���t�|�e����m?u��/{;��r\c}0tn�G�G���:4t�C��U�[�gݙV=Q�ی���Y�{~]Ƞ�4���:�g����L��%�/���-
�����c���t�k��i�T��t�0G=�;̾���O�s��x��t�h�����Z����"�5@6��ȷ�������KƲJ	��e�b$�L��t*f|�芉1��LdVߚ��U�������Ի �Vx(՚�:�Zj"�+�	;�(��:��5����W�g_ң�v��@��=������H��p�MM-��|�łԃ�ޮ�?&Ifܯ����@��Biڦ(ch���;���@��{ "C���aDéi�i�e�Ec>�xE���=�[�������F�
��ۊk�ȷ:���0�p����k�ͭ�y�d5�h���ό�ư%9�1 ��cN�j�w�������G���c��$]d+��m�רL#'H�t�r���(utm��K_�eյ��n]on���<gN�nV��D�����'E�"���J��D�qT�fHhe�J���z�t�I�����Kڮb
���v	�B|�;e���.��K�b՝�&�VӔһR���x�J��FT<���\��� ���E�x�B��l׾���On5�f���8�Eo���Nn��>R�)�'�܈X��^C�+-���E���goQj�v40|��x!(�"�"/�9�߮[^B�7����Ä���yn-��E���~n�ͯT�S!�Mb�޹݁�H=m��� h���Es��J�:.���z�FW��/�T��j8����}G��|��S�Oo���[k��7h���x�|�ٟ�IXu��^UR�P4X�ӳ����֪Q����nsE5��fx�O=%>��K��!�B�eؤ��µ��B8��gS=~��DY��D��T�Y1�x�O�'��o�=�� ���S�+��ռ���6����.�Bdjn� �ݘ �e	
���z:��-�;��ȵk��hj@C��Ϛ�&�~��q�Ǽô��
2�}���!���vG���t���0=Bx�|	
cF�d{���I��iEa�08R�]si�H������ f ��@/�E�@Q~zw�%��yA��&�7�>�,��OK9�θ?NX0���Ș�OJ�S��h⼺�r �,���,�9�O�
N��_�Y����%�QۼB��(@�&H���<�V-"OR���u��� rػ����՟����M��k��g����:H
��[;��x��j��Ҏt-��J���5]L�_��6�ǫm���z6��k!���.5����ʥR���S���#�4kwH���W�y������H�cE9U�D彪��0��u�`-&{8>�-�����ՋW���[lF"����[��U�B�xxԸ����l@���Sǳ(h2n��<م���Ç.v����<��U�_��lIRC��������7������W�HP�F��Lf�PC��va��\"zl�w�������uWGc����VR۬���"L�S���vS9rV���k�ԊO)BI�2k�#�ج�ӝ�ݘ b����E�� �i\��������*���F�)9��95y~B��l���u\�w�J>�%�p��]�>Wg�����;m�{���S��d(o�~���h��QMt�&��p/J���{Dzi�"��L���H����7��$\{3�g�I�?�f�\!�A 3��]����Lϵ�1ma�r��i�F�ɧ�����!z���J�S�	��=M<����] ���M:�z<��
�@�O��@�q�ba��+.�W���q^2IBHYU(����:+���d�6�9{�g���_��o5�s*�b�`'��	"�nf�r�	�����qD%G�K���o��0B#ej�%��2Τ6��}6�����+X0����w�@i���]��|`��a���5o��|^i��=����W���$@`u#�&���MFY� �������u.Ϫ�
9
��f��[>aS���Y��1 w��;�n�Z�%�T� Z�bوe��Q�5tN��Rt-3�.�BV�ITA�N�fQ����F�,İ�Z�����Ɛ�9t����v��Ѱ�q�U,{E1c1� �'��Z�K�|:jz� -��о���bش/�(j��r���r�Ʈ�1^N�3?7"��G�������K�����qL��������KS��pN�y2ӆ�zJ>�q[���Ɵ�F
�S�$�S.�:3�!-�y���IZ b\���ӑS�S� �B�6C���2��Z�JpR�����ʝ����Zg2��`8�w(A��c]�N"Ǚ2�(��U5:���n�2I���L��PNR�W��jBķ)3]t7�%����.����b 8�BVe]���ǤfF5UQ��?��y�]���!0rUp��C���u�?P����\�Jh�lft����(���|��v��E�&7�b����S��z$�<-��IA�6��{ӌ�;K	=�wu�O�#Ъ��bn|���p�a�-��i�1v�ူb��z�5��I�;�Yi8�Z��>����4>I6��.��o-���/�&m�9��������T_��E���t����c"n�Sx{�&#7����	�뜚�.��}0s�sG��`s�#�q���,����^�SU�L�`v�g���	%rz;;y�b�H�Jɗ��Qz��^f�x�=ޏg�m�py{#,p�|:'��t��_D�#�γ��@P��Ca��E�����}�$mtSI��1�E�h�\Qu�8�'�Mx}v�`�S���J@Ժc���`#>q��v�3����ǐ�O��
ĭ�Z�%�7����~&���^���f�۪�a�9u,j�����`�κN#�C�C�����2�*��j/A?a 8����"Ď.BT��=���Ē��y����TN05&LnF{A/\�,���K�ǒ�8�0��#�&��%����ᴛʷ̾\\
tN��l��%ȎK����IV6�S��\\�
m�oLGD� "�7%��q�%5O�]{�{H��mah��(��,���?��V���������tr��R(�֫��.ʓ�u^J��1�J���v���%��1C���e��dqR�r}�^����Lo��1B|�
�,��>�����^8Q�0��4��`�iT3�q[��D�p���%M.A�6R�9�k�� A������Z��x�*V��a��$~{�T�ڂn��.��ʃ*�'�9~�K��LM�0�:�U�w�N��[�	K�z�q����~�pǣ# Y�<e����_�߉��'d,e ���!���=�`�%�b���x!&�mxd�肩o, >��Ie����Z��y	$%�� ��8�P]=�Y��.G���dwK������fdo��1/���,9p�6y8�B3��ν��m��G#��@�!���2��$R���sc$�J|�-�(����>������y��~ڎ�z�k���P���2��Xq�w�E�<;{Ƙ�
�;�T����[�l_�r陃���ƴg��Q�۲\H><�RT���|�<������'�<�b��;ĳr*OA��̯�y�\{!�B���������S)���  P���$8Y��(��<���y�����l;���e���۷��7���:|�?tP�pEa�2�t�бd����ʭaޘ���;u-m�w���D�/�0���g�׆�����+�/���4���k��?�T�,��Ȧ�A�j�G�aHʔ�
��Vo�EpYD�j��zJV!{�7��ӵ�3z�>�+�2m8�R`i�̸���l�/B�3��@�ʃ�/�1�9�r_'��4��w�=�!9��� 0�`�����`��st�῕KtM��zk+v-��4Z	�l	я4 )[��k���mS� �	9�>Z�@4&:�{�֌O��B������e��(�'wR)�M���vè�����9ۨZ�U6	�^tVkϩ^���y�Y��_��~қ����:*L�$��6��h�aTM�ش�\��#�ŞS*����X0UU��#������ĩ�;etQ'� 	hƥo�t��qZZ�x�o�����~���!uf���Bi���[`�}o3j���g�!�O�Ӹ��X:�%魝�����w�K��ߕ�_�I[T/؀ģ+��zZ`3�ף;O��u-9eXfaAg,ņ�!���h*AW���Rs���ϙ�ǎ�;_��� ӏA����*T������I�>s��HF��k�����b�.�wAG=O�Ա�V�J/��۪^Y��䥼nY~�i g��!��X~؇��e�Q���F������¹:%",�!@�u_G�:!��S�V5�v�pE��_l�ɬf�k�*AB6���_��,WG��5�@��һ�Q?H9�MO���p \�B��|yҥO�)w.�a��mv*��7a`OS�"F���2]p��Aډ'j)��ϑn�?�s���J���΅X�?���T�*�l �^��+�]B�����rX7M;==��Y�������3.��u�Y��+����JI�JV;���o3�S`WŎ_�xq��2���7�Fл��� n���:݁�C+fe1�`�I�q���l���MС���������{I���:�l�7`,j��
���RÃA+�Ź޷��������b�=�v��$�L�"��bey�9F���bL1�1�����J++��C3罎E�W��flc��1��8C�c�ƭ暼�F�-��#m��7M�NLR�jJH�=��FD/�����)j����t���o�Ρ߼s�Coگ��`�	}��z6>uM�����uD�A& D�����w��ϗT�{y�(b�8�`�l��"[9�B�4(-'wn�QV2�����]�g&7�KwB��I���n�t�R^V�D��#����}�"ˮ�bg;��*���K�ucj�~���d͹Rd�&j��ʐ��i��ξ5�,5y\ғ��B_�D\dC��ɱ.
Z��z�/7�8C�#��*�͹ޘa�1����$[;n��d���2i��|cuOYv/�Ŝ׭ʫ�I�v�xb�Y��Q����:�Lx�]����	���S��=OP�K'H��	�­m���4(�3m����'P�S�ɕ'�I �4��zF1	U6"�y����-��T*7O���q��A��4]���f.�i��=��^��9^_x���~8����{JsX*�����j�wI>Nn�S&�$4���=�|]lGxl��A��34NUMRz:�\�a�jcd�E�ũC[l}DP־�����߱?B^��%�#���tdl�F����9%�rp'2�sXWwH�g����\%Y�p��)r6��(Fms-�&	�����o�Ɯ�$��y`���ԝo!�k��Z�&(Ec���C7�z��mK[�-��m��x����n1�P1���BHŮi�uI�O ���@.~R�ҿ�K��w�#��`ܠ&K��
.��j�|(i�aR'�U��W�SR�� �sa�j���p\�u`wsqQNY��βv��=��,��&S���Ⱥ>��)F�T4;�'i�i�a����]�#���t��Y ѳԟ��+�`.���q)�)�4"�@���\+w:s@��D�l����ge�'?^���g%��#���!�[Ae+����;�a�z�a2Em"��{��^���r��(�O��c�l
�`ӽ:����$X21��<G���+�^��U��'=2r3Y�tJ�?�E���l�(�smc���lZS��c�Nm�+��d~�		Xn{��D -�������X�u�8�[��Qt��P������N7F��ܚ�iպҷ@��Z�h����*��U��TT�MpHPi qaW��[p�}(ͷ������?=q�dmZHI�@�齛�:??�����L��ճw���s�t�o�~F��� $���S��_l"���ph�mqu���l��gݲ��E�m���".���V[�KI-�(��Z�%����O� &�f�鰟a�U��Ʃ�K��_�g���t���%�5����kp����wwwpp�����w��w����ڵ�S]��
�ص�������9?�u�7�@����y�#���w�l;x��!������L�Iݘ�B��/�B$��-��	�6u�oƩf �08�HTi�z7th����Ŀt�]|�@��ۜ������g^uNh|t-8���F�!)�Ni+.��X�:�A��ᇯ�wוu� >^R��j^��l�~"���x̸' ҁP7��?(���e�*��2L���M�濷�D�<Ԥg[:ak8
�y�Dr��q�!MS5����N4�����#�;��l��n�5��!%W�V�@�;_�>jN�Ĭ�	U>��1nZ�_!��T�_Ȭe#w�QQ:M^�p�sge�żg���		w�~��:��V�K��iiK1���a�B�}��4�_�� Be��9�B��6Oj6�e���������9ֳ�D�{��G+6<[��ئvzp���ғ҆/�7��婋S���2DCiGx=��$�QQF�AÊ�Z�<�!��I�d�����Dal����$+Ն���ҕ/����c����{���6HE�|�Bi(�,�3�R�'�[��ĺ))�V�ԩ?�A�Fss��L+Itj�����^�x"�fm�6���*$s�̋��~��qR�&��bi��d#��X�Y���V��}Sr��+��K�;��Zg_�ܾW��a�6�$S��Im��%(�J�z4 �h���S��h+��}w�E)x���%�ʡ*�l��*�2���V5i���^"R��{��M��"9���>d��1
o��
��s��&��1y||��eHm�mt,�1?/�`�;��ܷ��H�������w���>�ϙ���C��(V8x<"��j�>E<�Uu�A���7�d�����0W\��MY��ӑ!%<���]��H/4'G�Mzs�b1�,77N�d̓dg�K����=��LGc����������e�?����p�}��Kk����0%���8����3γ$�/E_3��MY������H��@��nV%/8��ݪm���Z�q~�5��`���V��v/I���-�����a�<�O�l���?]�B�"�4�폃�I�ؓ���DN��|��)���ʦ?����رc������{�����ss���uΣ�yW`�').E6����62���� ����������oBm'
�{���"<n��!�}�i�gY#�2�	�c�͸�6ZH'_F�a|5���+ŗֵ��Y��tN��i�M�.��Tmn͊����NE
�<~޿�d����p�
��x������<.v�wq5?4'��=��������O�݌@(�f��u�ZOHO_ٚ�l'^r�wܦ$��="���]&�7�
%H�l��P�ش��q��:0���.���`�vW�t����Z���J!b��ϙ)��0�ylIg�NXdkCmc�k7;�ܞ��hLfWh���ZF�t��b���K�*�js/z:�E�P���g���~IRx9�L��Ɛ�"�tG��<U���wJ�Fa�iw*n 4�)�|m�ǕW���x��P�Q��Ym4�g;�n�����{K���"l������N���%�>I_�(��'��yem�x";���8�7���e�4�!�	��o��0iLÎR81�p4N�����J��$���c�c�yPMpE	Z��E�/��Bw�c��1�d�ÐH�[;m�i
����qE�Y::�I �b��<�R���y�P�|���o���8�@W�||����|�G\$]pX��1\���M��FH�ԫ�tri�q�x�s|�#��:�#�\�����6��_̎��\��W��]��f�INb�.�gx��Bǟ������& \���HN)ǁނ,��X����&�X��N�cb�=�+<|-k^U���{S��R��M��gk��_EC�;�8.<����--/v}D����
���P��lF1�(��o�'pӋ���ȡ�r��j�p/�h�)�����m��X�z5�C�W˒�z�9���L�f!+&!��n[\�J_i�.?0�R(Nlދ�V�P�0��Rv�魞��L�=Q����Y��q\�g��%��u���NM����H��H�/��=%T��a�J��0���$i�'^w�謴�st�p(k��6LiL��9��i��d��7�k�C�!�;@��p9�q6M2��� �y.��|�55��*�Y��{�=��v��Sf-?o��K�mm��i'�q��;���u��������o�����|�o��5������W��8��H*����d��e5W�|����r]�2���]K��㙳�c��o�,�b*`je��R�{9f� �\JB�J��k^�}z˷�K�����f�]�cqcIITО���V�caxa!u+&W8���
��c�`��=�cA�(0Hw��uz�c���Qa�|R�>���UR�h��9�{x������J�����v��;���iH <�'g�\^=���\�X9�z�e�1�M1�C϶�Q٬�Lm�	'/�Yr�z<��d�V��c��e	�ɵ�S������YϠ_ѡ@G/NA ��D�t�@h*׾�-�I�*���R�*�tz~':�1��8��=��'f��Уg�{.��v�W�k��M�4��y׀bM,
݋�6O�z*CK�ґ�&.lcB>p�X�7Oq	�:m�E��c�+��QkwЪ�/x<zW���G�Y�'Q���}noK�F�,��]��ڽ��������� ȱ(��>�^��:�J�.� �X]�`���3���3�-�����.����`�������W�=O��&P�͖Ԅ����-�\��Mx޳�y~�v�f���5͎��2�~O:͏j��E"�̰��[�S��/Qς+˗T�)z��f�(��-���X�$��9u[�J���y Tp��S�W!�k�ú�fP'���둃�Y~���˔��Y�_���k��m�kMߢY��-�ǂoPb��'=t	���ax��0�ŕB�����2p�詁r!�Eͫ�,yZ�i���ި2�����7�1�{�%�(�M�����L8˴l;\��潩�o��<t���
��ś1�9�B]�S�u���堯}S���m�Я��v��9��H����Y�W�-j 35�}L���4�����tޛ�'��^yZ7.�Z�L��`���x�V����<a%҇A��'�C.�'$ ����y���tZ��A{�2�K�^�"�WU��!���������J��.�:����`�)4�7��b���_ ��<��ڗB�zʥ;�|Ȱ`��df�&5�TU�uW�XzGDm�#	g���zx6�wɚ_�g���υ"�lsg�NL�Z�Q�)�k5�4Ȋ�BѾd�g��;oy1?�t)v�>���3hpC�]0���q���p'��4�U1��Ֆ�D�&�5�H"�A��:Z7��X��e���ZM��&�7��Éav͖�-��%�{C�|0}�$��g�oUY�z�avk5���܋����_qU���T���8�5���u�W$_��H����U�7n��|Wt� /�������A�T�����_ہ�sb����D�e5=���qgG��j��ͷIJ��W �s���Ҙ� @����$�.WE4ۈJvAj���&�z�P��a��b��G����(j��E��nq�=V����x�]g�7�|c��F.�&����j�x��P��$k��-OL���Ӿ/M�����Qd�a!��H�8.�#L��R���U8�1D�֚,�Շ] �u�ֺ����h��Q�<�x�\2��~���н���� &�,��QY�s�A]v_o���n�dL�֪P|{-2tKg��R���ؒ���Q�����T\ЛẞDغz��/A)�u�L�����[We�l��I4����e�|s�4��"��u �Dl�\��]i��<�a���w���¾���w*�Y��4�x(�V� �Ʋ4ׅ��q�*Z�z�u4��Fâ�Rhn��Y�<	`~ˌ���i�#�ab���Ö�V�⎦�[�+�w�7%I|�0����g��X^�Mw�� ]FX�qmir�m��:4*��C�����[�lϒz�������$��蘘	h�_�f�Z�I#�8Rc�L��, �9q�a���+�0:Q$�lܦf�:Y���@��LՐ���j�\0w����%���(Tc���l�VY��(�l���7���jq5eh���.!��}���x˗���!-�]G�¹ll-��$b�I[�gp��r���k�M�޵��#�i�_��a0?9"�<PZ���¸ @����j����k���c�T�g�(7j��vK�zo)(\H��)���)��,�*
yeq��g_�����d��8��	,Ӗ�&7g^��#/�Z�u;���/'j���i�)��|b[/��Z�({�O�E���T�j�iD����MF'3��}�)r8��d��M>�OO��4��ŪP���` �R� ����o�����p�N�Q|����͝-�F~�!@���U�9�;;t�/˛Lt[��{��P��*�#��Sy����i\�M��lyLwmƱO�'��C$�i˧EN�ِ��U.<���;��!�-mPP��&f5#o��[���_����o(�ͅ�GwL 0�Q*j��cJ滫�)%��;f���J���>��ܸ�B>�٢;����+�@�՚K?�:tc;��D��g1���	����v1�
�O8���v��ԦO�l�"���p�Q�KXIip�Е˾�@�@H�k���J{۰K�x����'nUrBu�Ձl/څW51��Ծ/7-�m��Y7�F�C��m�r΀Y#��Z
���JRGe�I�0nC��E��8�WO�v�O�"��{�lo͸��2��������0�4�#�����Tvv���uZ��<oh��DtEHd�΃�uX膭m�	dC��K�a)\4u�v�鯲q��e��_/�k-�ߑ�_3���Z�*��!0069O5��t�%]e��f�����>@d7�A�Q���<��cg�rV2��O�����;�a���#4�Si���c�J��}��'�#{��
d�K��$�s#�朷�#��.�I:�}	��	4�;,:W�m���Q�����A��Ky��
%t�fa�a�RJ�L��8�<ӯ��D:�3�{������<W"�4�	{�ge\5V�O����|ګ�_���Q���5��`�e���_���L��;���"g�]j���|&�	�:�<����/ԭ�0������<�}��F���Jl��)��V�@���k��@g��U�sɲ`��w]�Jx�k"|˿��&�6kMb�M�Xa�J2S*�E����nM2��B��rOpS���
۝�����ң�t�:���>;�*�@��@���*�S��XD�d�?��~*��i�]����xm�Gh��0	B�R���>�2qt����]4/J�k�o6�/D>_���Sg{#$�#��)��
���cf�:�Y&�SKwjNTI8�F����im쵉
���ok�@'��k�/�{kF9��4ՠ8<k qҘ.�F��?DXF!Qڵ�w������6�]�(�GG%�f>t0c���L?��&1��6���L�t��k���af�H���<)�Kh0�䌸��ÚS�ڬ�z�"�z�A8��o�������	z���U�Im�$Hކ�&�o�e��=���c��w?-���Fr�٬�C��;�v�U�j�L�_��ާ`�t��զ�_���>R�}����"�����z�.��I�p�s�B+�k�,�2�-��y��3��`/�� ���V̈́�7�a�tw��Ig��q�CW�©���׫�X�Ix�-+�w�	�7��M��cu�.ՙ]�������g�����ݼ�_�vV��/��[��H��R���[8���6�o�d���:S�`g�#��އ�98����U��@�2�!�[�����D��ω
*q�2k��������N����S�"�J�`xdM*\8�,P"�K�?�T�a���h�<m�l�� /�,�H��`T�ٯJ��Q�����3��6����!M�f[����]ޜS�t��{�ޮ�$�H��w8�n��imU�k�.��c�A�Y���|� ���:�$�I6+��p��'t���#̻ ��ᐳ�����8P\!��Vȱ�T�D,j�rv?Z��u�D������{��s�eِ��[�i2UF4��ɯ��p#�y���x3k���A�����!M�V	Ք3�Y*�O@~֭{m+ ��7-/F���N������P>,�F�.�u8����8�~ť��8�6�a�T��[(q�r�ׁ�P�T9��-c�������L�N���� ��G+�&��?O�1�$���y���-v4�[ˑA}5�t�H�Z]ʹ- UUt�O���SJ5-�A�W�3
-�F�l]�/�l����-�X�#D<ovX@C�
�b�Ml�����^B/��T��!bm%���hh\X�w��**�Ѳ���Ƿ���
(��Z6I��l�F���d���/�7�R�=A:��&D��ٌ�EA��<H�F�Xiy7�"�(rEڼ�WU����+�{;��6��vyIqh8�y�>�a_X���G]J��>��kW>J�� ��ߘ�J��
~�u`	���8������QyB"�d�s�ka�S`�ئz�sL����t���'�|A�Q-���Bv�tZ�)u��h����m��B�h�&w�E.��QX�f]�g>�j��?t���4Jx�>+�>��~��ͮ�����rZ�h#>N)8*�\xh#:ݰ�5��ϐ���"�t�ˋ�a��GV|�,E�T��z���n��.Dؤ�i��9�3�*�]{��.̝F.�e�|�������!9/��^/9���:KC:�>��ܸ5!?�E����D���E��������=: �bt��GԊѱ�e�"gd��ۍB4"q�.}�3�Ș��W�}�Kdjr!	�ƅ���T�#����ҧw]�4�ԥM��M�v�B�@i�o6����
��D�y�����v^ ���A�g�S��v�q&��}�$�7b��VT�������]ioxQI"�{;��c*����*qN�F���o�(�p��Q��Rnj�V��j���,�4��0�L���>MB){ ������\�Gx��@'Yџ:�g���A$h�����$7�\�h�1X�H�G�7<&�_��˟�mf�mG���n�np�W���(�8�d��C�kU���Ub|�z���X��}d�5�Q�Y�~���隉8 F�.��%b;�b�E�q#���Ӊ���S�T��e�HߟƆ�dsb���e�B[�]�������9+�yaY�-'�#s�Վ
�;����U8Fk{�'�FS��S��*þ�a���zȓw3�c���vy.a�}�V�#�Ki�6��bZx�\X�b}�-$������ ~(f���!8|[����I����=QX����8&��!��٪��?T�0�}]̆�C���݃�b1Nlϵ_�+N���;���bq�N�Է#T��u��_�)&:�K�$�����d��.����A�`Vm|~p��0˾^�D�R��3A��;TW~��1��}�N��#E��W���+��0������rÀ$�n欵,���B�1���|��'`��h��t��(덹�ġ\-�~�����E�)oM�k,!a

v���Bg&C:]d��-,���9W�>B��y�E��ww	�g��5;D��������rBq(�N�ж�;C�<�%f�>R�⷏Ӡ$����?��y�6Rbj�v�7+M����l���	��v��"m%`�/,�C�b��h
������,�z�~V�-:�62� _yO~3��B
ٜ�^�|��"[�~fj:���'����-��&�%��!1j���3:�,x�z(С���`;�w(;��^�4�}h��?EG�g�����c��a���41ך�a]���C���!b+��n.?�f�9&E�fÙ�w��4}��C.f�aP�M�k����Gء�P2Y��r7tO*WH���������G��dP���:��k�|^1@JlcU~��㭒Ge�q�b��\<۹�J�Dʌ��M�0�o_	%��`��^�q\��G�+����ޭ2V<�,���-�����9Sh�C4%�[���M��譸�V�L�{�4�3����A�>�����7���g�K��#&���P�qyjc-ݘm*�/+^�Ap��cDD�E��V#jUI����ex�=����8�YÝx2��SzB��C���T+�L�$Fd�T⫸D��e��ɲo�d����^��k<!����5���F�h�%p�$
�LN8�ﱻ��y������g��)}WڰU�պZ�n�Ǧ=]��""谱���^��rSr��z�Jׅ�5[��=��d���O�X�����aMk���6./��=�w�n5�m���M?f�F���z���Wt�A���,��6�u���bgr&�9���x�/DP��f4�zau;�C��ܵ�%CS�W�-��N	�9���S>i�|���ǥ��9��B�[�پv{I�@���W���S��_���[�0'\�$+"b�Dr�a���&ʼ?����47dn������	J#���L��9����9��{�+�$�I: ��;X�q��hSH2_�r#�ȿ���<�n?�<����Y�f�@�]���w�G����t���:7pn����g��.��p�L���o����a�9��LQ��-շL�J���`�}�ܨ۴ut-����Ka���u�x���O�Zx�����e��ux�a8�͒d�[â�o��=nŧ�(	�����K@Z'��F\�%��8��/.ŃH�߻1�dg��)���3C[Lit�ۛ���P�r�`������,7d�����%�1dSI�����=D��!7�pS��"
�[v��~��W�?*�(���5��0u:S8�i�kA��b�`�W�A�|O��Ɣ�2�ɞ׃;�ͩ�b����2<��~�ӐX�(5�7
�mK������6�x����҆aZ��R>�k5�y�#���3�y��S����[I�jO�@�P6Zz�����6���bX�#���\u�F?0�_�Z?���+��(�\�N0{ó(��J�#zW��h"���x�1�Hq���c'���VE�;&�E-ز�(j��{=�_*rk� Q�',ii���� T��3O>B�
b7�h��F�����͌����]rX��gs�e��÷��:�u&[P�^�<�ȓ�Uiue>26^��V�g��"
j:cru�i_q�L�B�TX�"㶂����u��hT;b���_��S[Ҷ��jG餴މ=�(�4'o���w��B6ɢ�᱗��)i����-��a�D����%�f�©_w�i$����(%]���=�6�txu���↞<����&�.:tc�|&����Ƕ�P�F+�k�(<Z�����yP���%�`Xtks�9����X�b�z(qcV8O5Y�
W$���k<�l�3�db�0��>�1����r��p�Ϳo��TӃ��ψ�oJ-<�k{�zJ}�|��e`��{���Ĉ�wNƎ��͔2��,D�-�詉�]�^
_+�w�ѩA���`���#"EH�[��"C���h�Щ[�Y�-�Zs�+ncC�(СkG`�%�l�/����;�����ݯɉ;�gF=� n$p
�e]���/�����kk�G_�
��Y��ݬYPk��֬���E!�r�Y��&�p��9����A5��Z�I�,Em���o��H}ti?d�^�F�)��5�N��㪖������ -2*{G��ƣ�x�a�����V�i~%���1�:P���#�3'�+�k��78��:�H�����Ґ�-*��iK�����2�:}W">���^�_T�+�O�J[�wu2��
0�S�P�ɭŧfg_2���qM�l���~G��������Կ�?>��$cC�������%^�r����KD(9X�hs�~�7��� �o��WX�[��ZF�����qj�&�h�C���ޯ���7���oh�I$N�-��Š`�­�^�(4�;�V�19������C��Y������Vq�1���u�w�Z*o�t���˪d.���TW���R4ۨP�rŬ#�wP��x/�z�x��[���>��Zd����Y�f��	�3`��JO�����.8�(�,P�`�$�������B��4��R[K�q���jǙ4#C�zF���P ��� �~�G�|h�����<S$�+��.�d/��:Ô��()�u	�$��´dz�� #g���)�rD"���|�e>� �1���o�"�Xǹ74�n����j*P�b�a6BEg]\}���J�++I�����1�p�+�o�T�#|���9����%�8�
��	Gе�F	5�z�H�o}�4$.�Aq�09qn0$���E�#�!�+�K6ʔ�]���jJ:�P���ژ���eNJ�4V��?��VG̞�Voۍ��Q	��mE�Vl6 �@�
aԥ)J �x̀�f%Uʹ�]㹗ҫ�X�������r�*w�g^���)u�ݤy�~{<#m����D`�U�4�������Z'-�J��9���ً�>��`����7Ξ��Λ`1��1y������=,~�h�;�,�$���.DI��<���t��3峥.�i^�)3�ށ7M����ܶ�y_!�M	K/n�J���ז�@d��&uR���{��x(�5�a1�7Bn�ݭ3�C��p�_qY`��i���6�8�xIɷ��϶=M~`#������ kx�;�h_��KG�)����lb����[�Nq_�<��*����<�0HB*]�k�2	���Zl����M�m�!yOEz�;	�g�g���dxd��{G����_�TQ�c�+9��"e;:1�D5���2b���A`�d:ܔ/,��B�qw�P.},���8>�͎m�jP��9�W�����ZA��aU�BJyu���3��r��g̑�_��k�{�5]��̇mW���ɱ��M���!;����+��	��\8�?���4�#�k�c�ɫ78���9��� ��ǙԡP�:���ڟS�E�
|�ň� ����J�Ae+�b1��rh�)�i	���v̊[�$�©64C���ڏ�o�Q��%,?��.�T��D䶕��q��m��YH
)�˲C���&�FF��7�P�O�WF�3�/��'�4Ŏ�j��^Qp��8����\��zc�j}wkj��4���8�l@������)���͟`i���w��cm��-�ײ�QU>������W�K��4�j��k�^7<��cݴ�	�tf�q����U���9�(#y?#������R�%LҲ;��V�	r~;N�y.p٣� BƋ�l����J˘�۟���5�8�b���e]���K�uCd�1�ab��s�KZ��vC�+S�_����1O�?�)�n��Q����F�;�舭g{(mk�I�z�n��|��ަ[gq-��o�3S�_5����c+�1�^�#���H��6[|�Eً�P��c�V+<j#���6��O��|�s�n�z���4K�����Q�֙32�Z"�e�E�N�a��v8�q����c�wN:���Ɋ�Ř���F���ef�7Jl�����sen�wY ��a�7\Ra�s	�s��D D'�4�m7����
�ybҐ�L�X�����x�7����Ҭ�l�Z��kW�^��<lFW�:�G��̦J�#��
Q�m�M��O������A�t�o���q�G�756� .��b��S�$+J���!wɓdbc�SU�)���q�L��/�WAo�L9��^,�$�{����V;9m�����-qv���Q���W���y��#,�$ScC\
�U�7LN8 E�!�4�Yĩ�`��M����G�Ln�ۘx���0FW)��Mcŷ�����Y��8�`�<�Gkk������cP�k� J<�	�%���_�~:�?���w�[=(u��L2D6K��Z�N�&�z)�gL絩H��#˿�|�t�X��j0/�ГO�7�Ҵ�Y�\���]����M���ƆG�։�a��U�F\��X���T�܋a�Mc�w@X��p�E��'d����-W��m���Y�f����k�)7;>I�� UUl��;e��1�9I��5�."����ȫ�|�[��:�
%�Y���ے6���� ����~6ѕ����-�q1V�Y�RB���)��_�c
�"��E�t �f�������*��D�X�Q$^D୻UV�.�������.}����3O���t����#.�����2g2��r�t�:��,�Z*݅���C�`�łjz��H���-P��ܷ9�Ұ��Y����[�_cB?���D��40}���8+�5�i�	�/vU�Ü>:r�m`�������4��T=����6�f�*oX� nX��qLb��������&�?��O������1�@p�hy36�z�!\<��*�-r?����$��E��s���M&r�3���R
���*'�W��'�+`��`?Ѝ�8�U���/rpD�6�K�¡�Nl�wr6����6}�ަ���>����1�A5���b�?ouqY�2Q"q:j���l�Q�'x\\T�ȃ�~���7�&��<�]º��C���a��ط�0����~Ye��E�K��u#l���>lLi 1�s���'F�]6qs�T�G��D�@e"�� �R<�̳��#�g��.A�����I|��=���"��`����,��a|��В[���|y�*v_�鑡�'��q����k�z�1�����q��^�V�Y�=0F2���{��!�H,u]i6��dS[B�e8���ڀs��s���%@�(?ȔG��X�wj�<�ogɸ%�׹j����]n��QR���lG����M::�|�d�Ӧ4���8��s�GF  ���8�0���y�')�����E�L�@$ҏ3�Ւ�M��v\r�����;7�c[Pa����٫E��XNB��F����|KwF�u*����>�l-O4Y�틎�'Q���aѳ<�Շ֕|v1��G�i����1(w%7)���]��n��%�%�܀�qeR��4Ӆ�Du�4�z�J=�|=,����<��/2C��^��2Sל�%հbMyJ*��m�ʆ�q�m�0DnMNT��HR��� Y���	0�zӳ��?�a��23pa��(:�K��И��1O�ɻW
����������Iy^U�L�9JAs-!X��/���#��d���]Ͱ:GV��K�ACSϨ�ea[�VR�59���P&2�j/S�'��9�S�dԛ�.�>JZ�7�M�s�+�d)�x]7\^�)eȲݱA���G�6��(r\�"r�<���W:|�5-|hԘ��1�b�
{��ߵ������7O)��vMΆ�7��q����z�}�J`�I�d�Gtl�?�!�6><��������E��N�ʗ���6�T� �]�L]�E��r��&�BC��ME1O17�+ѦP��<�������;�م�p'��Oђ� �"����`��-ҟ�Z<;F��-�+�Jr���/�:\�NXj�^`���a}v�F��7fBԊ�j���!�cx�}N��%c�P�R��Sv��Ч��'V��Goͷ�(g��ߢ�w;�ܠ�<j?��O��&��$�(cZ3��J-P^UcĒ��dlc-(霰{H�Z�h�6g�O����o�h�]7´Z	b�q�\
�>HI����8�{��C�Aυw�er3��w[���.�|4F�VD4,~5�i��H%T3
e����JA7�f!-��n���-�҇���X]M&?oB��7y؞.3f�U-{�U'�G�<��c&$&&�����Q/�f_G��C"݆�|3,i�rJ��pX����esӬ#Q�PQ�f��ůyt��W0ov�7��zx��d�t������y�/�[��h
u���&.NKRD�f4�S�[+�6�?Ac��#��>b�+ ���]
q�`We�.rf"śj�,�t�x<���+�e�����}�'�Ǌ�D�_�~�S�G,��V�[5�l����Ai�Bt	O�i�A�N��Y��MQ�>��䛽��_��MQ.�������\�Šv�����T��Hw��D�B������үJc��u&���vKH�Ҋk���0)��Ntw�'Nʗ���������p�w��[~��L=��bG}h��/��o�Z�'F7����ȁ�8� 8���s:6��h�����>|2k>K&b�qb���b��z�w+�[�<�4��&z�ei(<L�'GS�y�D�ǲ),d�����̑Y>]�9	^Q�R��	�
 �p�����堊Po�%w�k52)y8��YIIV�J�?r���^�?х��6&�T���ڽ���)�6] �G�ˁ�M��Ik;�t�O��%r
��x���2�x�5k�Smq!\����eH�.�9�韱� Î�ts�Y�+e5�{i� �j�������;#&��o7C���r-71�̙2���W���<hJ9��?�_SE~��U,mҸ��!�#�Ҹe���t�L�X�B��j���}����Z�j�L�c^V{m ZsjZd��:��m�Q麗q��M������7����
����\�a'�>K��.��U���LiS'ұTT�<��7�E�Տ��w�7_&3W�[ '�y�*﬇��}3���ܷߥH���eh*��l��n����x
��v���yᤐXm{�!��w	���F�PV~��F*]	:�Dv�P����9_�z�:ӿ&�l+�z�@*���3@�a5�<ۑ�kE!��V|�����wƜ?�X'u�C������L������fr)﷜$��@~8��k���i17���;��)S�y���E���lE$eFVÜ��2yS"�9��]A�jLN/D��3�%]��3B*M._��fͪ�C��i�mcN�� \�H�,�����w[�9���;b��Xfx��&7�}޾����K��o����H�.y�|��o����?#lُ�,b6c�d#��W�8orw�n���ޛ}>�워���rӗ��xp)��M���z�i�����XУL�/N�,�OMB��Fx]SN� �{�����ڥ}��PN��lY�%��K7�^)9D��"#�z]ǯP������3�?G# ���X?�V��řO\�Y&�=��-�Gxnя��n��%N��_V.�[Y�\�R�~��<|�	����D֥�e�n��$�w�x#Y)��&�'���@q��KD�L���c�Gp����\�Y�λ�͘���e��%T��z��Z���K�����D��%_	Xם�fe����?@�S��2�Le��K6L"��
�<㗅���)p6�G�F#!{D�ůX��	ݍ���˦I�����.{�ds�1-��:^�u���+4{�9XlX|v�z�}�5�k�H����s�@�.�ȠJ]t+�H}�v�Vݠ��|���Sٜ͛3�b}ׁO�̾���"�L%h>�%�-�K��������!`Qs[ӏ4����k�9�E1���EX绚�Z�N!k��+{;��qy.�^!������;�]�Q~E@��/���8��&��z�uI�a�f][%v��;��5�B��^ *��#�a��?'�x��'d�gg.D���=gz���u�T�c�����Bv#篝�������IR������? NRK%æ�����3�I�rJ�"r���/�#��8�9As�������'�~�cA�vs��<	��i!V\ݛ?R;i�3�n�r�ا�R����2	PĆ��z�/��sXh ����x*��`rf��}�����y3�5� �`�>=v��N4�W]W�bf0:E>�S��"��bNUP4�����,9����Ug��ڶ�:��Je���&M)} ǄQ"�<�YO��Kr?Y�[P��7���M'
r�@�<v�X�����K�b	���]
�=/�R�Rk�V�7T;��,s�q�������t��U	M ;h��x�#��)%*��\'9�MFI��^8��i��t��<���"ω~��OY��e�n$3��9�f$L�KlY��6W�^W��������fؚ?�hM� ����R��
0��� �B0�z��U��yɁB��e� ɵ�����\l�l�,Z��׻F�&`:ڥʥd]��5Ro��и�b"��s�W2�����?�࿑�#u� �������wV�(/�=�"QX=�@�����;��L<�V&V����͓���{Ğ���O�s�h��VQ�.$M������cp�7���J�� R��}����a��'ߚn�G��V�R�����~u���l$����k����Nav<q�|�kx�qz�T��Z��6��](.�x�b�������%�w���Z܃(R�w�(�������vw����gof��� i�6>Ȗ0��gp/��]5|��oh�.�n�H���G��)0),*�v��RR�<GewL.��4|ղ(�4�[��'!j":���_�$糤ۨn=�O��dig���[�6�d�-W:�8�֧��Y�ݽ��ݝL��8��u��G��vW��6t��_R�1�� 8�-d�?���9)�3-Cq�-���k�U�������̀1��+ORG~oSw�J�Y�O�����V�X)t�rSM��nW�mN5g�Aw������&^e2�z�"�3�޻Jy��}ހ0*�dK���o����Y�*�|����>n����A�f|k]U��q�R���Kv��D Y��#�%���(B����}� Ϝ!o�4&�l�|2z	;0�v��왼~��(-oI�5N�6��i����dD��cH�}���D�)n��H����#�$)[h!�����>���3n#e@b"��h=��� ���=��o�h�v#��q��ÿ��_2�3h���	�*�c�pb1�<a�79�O�l�*(7�Xgv���6�!�G=�U5�3��Z�0��a�.}�n���(�X�D�o�`F�׊ù���G���Am[�Ӧ[Q��G1����5��d�[���ܫ{b�ӌ��������=�,d�9�Ŋ�'2.���b��
%O�y�w�w��2��9>�7�]g�Z�~��w��	'Ū�bB�h_.��"��^��c�x�H'
S�8��O���G����z���b�ՠȁ��Ģ O�4¤��EEma���AP`��PA��N�Po�"��V�[�:�/Ɏݹ�<}:ȸ1�0�^k�����ˑߵ � y�2{�����*�c�!-"���j���8�r�߬Yv�ܥi��V/7#��g�w�e{;��^;v���W�X��,غ��[�3�K�d]���׮�3��cD�- �,i�3��OX2���9gS�9<ޜ��z� �r���S�.d�Y��^�oj+{�}}O��I�s��+?uȑ�y����k!��JS����FO�zzĺ<�]�P(lo����*H�tniޞ����s���J an�]�ImSn�ˀ|aA~S�)��l&�R�H��#oӳ��V���3lv�|��LpΔÆ��3����G�S��?d�"dް�5q$eaм9�ߌ;��d����[�b��cm@��[�x��
��E���3}Z��}�L(��ν�$����OP�˳����!t�f��``��iU=h�.�uJB���(�]Bm��Aα)��?������$���tG���j�j,F����<��9�\�v�ۤ/Tz�<�A�Lt;���U�����#i�؃1�Q�Ϣ���>G�����ُC�b=@���Nj�_'�I2@����v�n��Qs-�P1����Uip5o���-�>����5?*)b� �Ç���`��`�����@3����9�ͦ@��:�9��@�zi0Z��x�n��kN���{zb�d�]�cS����"c��[#+X��R�c�5���4I��ף���R��qAN7*2��}���dף�'\4���9��^JR�Ru�©��v]zw�R���p ���*�*�U>]�Lo�c�/g�1i��~X2��6ugɀE�P�{�,��j�Kp����C6�[��\ܜ��B��M.g惇[��J��1��-z�X�������3�8�ki[�f!�]��<
� #�܋�+�3U[[O �@�z��,U�y�g��PL���l����q���I�MUT������m(���F�.��D1���e�͛�M��x��	�[Ԣj�Ք���@�4<s0z���ݾ��q�4���=Q�$��(����s�M�ө��v9" Êͪٹъ����!9�4fmF�W+�"}�|ʛɡ�26�$Xy=Ej5
x���&5��値�+��7��\�y
�%,/5R���dh ���)`�"�:BJ�ҡ̦yFť�\��7՟ �4/׽������ԚJrf2�P:�cx�v�fo"�D�0�N��
�vW�e/d�ٻE��%#h��\�d�Ts�R�k�����Ƒ�"������<���r]5���r��Nh�$d��C��˴�����#�d��E��{?Ӿ���c]�++�aݘ��@�AZ��{��d�nx�,38���~@N*vu��͵��ի{G}8�W�+���&V}/�W�[�M�$�t��ۻ��S�)#	8Ƈ�g��%o(
��	~�E�:<t�c$Ot��$a��A!.*���F��iU��:��w��D+��o�o|��On׆���Ƈ�K��I��y�_vT��W�^0�I�a�������~\q/��\2�`��0M��y��%�ST��7�5�kH6���ӽ��P�ub��]�6�4�w��[=�؜�	p�p4� *!���`:�Ĝ uKպ\\Eed�P��A���ڱ-:G��P�~8!GJP��> [�ه��߭C�]%n�tgB�8��q��j�C=R
3�0�C�d;����,��-V6ϙ��	&�CJ<	~�5�^6)��CjCE��m�a�����O�Q:�����r��b���g����znD>�P�X�X�D���X������w$-ó�zË��;�o���TM��<pL����+�-%��k�=�W�p�hD�p�<�;���d����
M��*\d�]�P�J�Ӧ��r2�0���\C׷�{P��1����9��}e�֮b!9�<�Y�7��؁8z�z��|M�*hr��tB�� Z	%S��1����Pπ�*ܪ���N��'{���#^֙Ns@,�	�3^�{�qP���,Y�ɻx* ��JC� KѵK�
cG֊<=���n�ػ���G/�=l�
�mAmf���=Y�P�������ܒ���^TE���@냅�fn=Ju��F+�{�k�D���)L���T ������o
��GR�%��Q�����y��]c�%v�+h!Mt��CZfXϖ�]�Fu�WU��h��B1��ӂu£�E뼇u����㎷^�s�3ޕ�Ӡ�?u�8><Js�M�ܾ|�t���S�B90ËV�%��;Zjq.�w��d��v��2��(�rW����͌����5S�;������^/�[�̯d��Qd�k���T���<;J���Y����ѷ��_-���3�T_���84۶`�� G�r��j!ӝ/����Y`��|}f	�F����-ybm�&׭���,��ɕ�n�!㪛 w֬�������J��:2S��]h
w����.���c�����ji_Z	_��>|����we>JF��-�b�xbt?
�>3i[����R���pnt�L��u���%�?F������=���k~�ܱ2Fc�}��4B��P���4�,R�q���7Gea�ꊱaG�7b�p�DLژ:�6$@��.�����x�y�_K�^b�v#!��j�p�b��i��t8d�w�JNe0����5KI��*���h��O��T�%'YE�y>�;�v`�<��ф��óg�T16z��b�Vr��%yXf�Z0投:mB�q�(��$bq(����7؆�t����*����T:M
�}��'l~��nabP(�q�kk�f�1P&��t�I�B!?��u�PFޓ)�<��A��Y�j?GH���qk}#���;ĔR�����-h����(hE(��Cq�0�% ^����k�U�.�KF�1�a���l��v����&��p]N�JLtk��͜�ke:����h��݆"��b+�A����%~v_�g�����sam]D.`����H�l���6�j�s�{�k��w)��)�j����<��Ļ��^x88e���G ��(�=�"���a<�%�>K�ڞ#�Tk�����|}a�A92�=8��ڥ��|D�Q	�T�J�\��`�����a>r��aװQ��\���ؼ����M���ctޡR~3L�H����K�v��G��F�x�o5)꨼��9�/���(�Ѻ&��5V~y��~*��yQ�pZ��;|������Q�/-��� �x�Ф��*��?�J�jo����H�#y��d�G�������s��}qNI���-�f�~�t5F}��� �d�P���n���j����$��㗴@����;��9�i�=y<Ge\��-�+��Ōљ�4w��0��L��0��n%"D:�N;b_����N���a�M�u�h�/X��u��(C}(���>V�7�o����n�#�Á5ۓ��-3R�j�����u[�����-ύ�R.��}�I�V�͚q��e���{���O�\�m���tS¯RT���Rw�;����h��uG��Y��
OY�?^w�\�6�Y�V����:"K�D�L/PP3Ӽ�&�ɚwX5}uqsgW���4�LRIt�꧹�q�/�P��q���y��Qk��ap7�zͻ�o�v�Z� �� ������c�0gA5["�S,"�_���p;�������}�[7�d��S����wxr���ɑ�ɜ����l�t�q�(,�*���E2���~\�%��?+O��sp�t1����\�2�G%����N6��\�L/"�MS�e�ඨ2�<����k���S��㰤�׈JG:����A����"$#�3rC�!K�*��bs1�ۑf�!x0��w5E%��"Ёkj���C�#Z��wsÖf�Nb�����y��9�P���O,���99])��߸��	��eJM�%"����ҞG�/&�ΪGb�_�B����&�ْO�O�Kː5�����*}S������^Az���o[ <�P�NRU+·�B���� ��QA ����񐖸�7���w�_`T�=%�B�ш��ɫ�Q�n۲2������#��0S�}-���&@t����Q���$��C��:}��%s+�7i�U��2@5�M�#	彼�ثϻk(��&h,C�j�O�n�p��K���v>��d3��Ʃ9�@�sB`?�#���/����\��7��h�������h�D%����yl�gi%׾����Q� -'QO�\�A1Q�a��D$�8��ڈ��8.�ز�� Eq�P����>$�D�*��=�.2���oM�vwx?�/7wA��yda�Ǫ���P��Y����[�����5\�@�$��0�Fͥ�9����l�^\MOw�}2�驞>YeY9Ƶ�)�Ѵ�zGZˉ��/�v�'N]S)rz�u}�<����Xs{�\ ��,<�8{	�_1��b�s��q�mc#�Qd��a��R�|h�慢�FBr׿8����\���v��o�|�t�����͏m��n����9c*6J��	��g/Gv�cZ�о�J`�]Yж=����[��T������w�RZ$}���l�T�|@���{��^�2�d��F��%t��{Z���R�г�.��1ֱH���ݡHi4�S!*���f��$'?��d��L��_i�B�on]7T�X��Zc*��m�k�h�u
9� ��-C�QI*�	�φv�N����z����p�O�C�W��0?�E��vc~p���b�CJ�#aZ�k�Is�Χ �� ���B�p���?���Sr[�xb�;6�y�T~j�h
iY
��N>o(���cjlg������a���BW�Ţ�����T�cVx���� 9�:_��TU]�Vu!�a��7����Z4������,�y�b~��`�R[�D��L�A�P9�����[Z��$@V�n��k"�>+ú-Q��ɛ,�����u���M�Dv1uv�:�� �TR8�.B�>c������N�X��b�T�n�1238�{�-$a�ē�6���j�(����H~�δ�9��)���m��.���q�2O�	E��ZD�� �/
���BВ���l���%��0�)V�\[ua���q�BEM#9H\\5;��1)\���'j/���~��\�a�5��ۯ��
�:#���?ӾC^1y_j<Mj�/�Ќ�.��h	C%�k 	��$���10�u˳aݩ0��\ �>Z��.EB���I/������������QJ��� �Aa��m�-�\��6oҊ�IrM��8-Schn����z��G�/ɮ������ᷞOZPd���}�HB�A������A=`�PG3�'���f��0�H���|b�����m|衪"����V�UA������{��]��3����"�˄�R�8Y�������C��#�h�BB�ba�8$���@UE�4ZQ�w.�e�����'vQW ��yd䃝��{l��C� '��5���@3���!o>��V���Xd��v�Ĩ�-T���2�U�p��D�?�]�Z
���w6� T뗟Q W�;D�������m�75�/�BSo::e��X�/x��F�4�,
X櫫���|�����I�*����S�O�,|Y�-������:��d�]`~��J�M��:A���T��(��m�3J����9S�?��A��F����!(|��G�h�����{��&b�,A��;L$�G�oD���.W�5=\��0y���Vi{�A@ڻ��`��V��dL8;g/��Y&�4?r�e:�9^�m�6����x�&$�4��&�O�o�%8<m��L"d4ȵ�����E?���ٿ?�xs�&�b��t�̾��]���j,A�}D'2����D�h?�9�*�?Sbg����U8:��Nf`(��xV���9xu`��؞��o^)D�N�NL�`��}	�!FFH�M��+un���h@	�M��D5͒��-c/��H�Ȁ:2���'��(��Ҁ�.�r���C$]����Z�P�B
e��/�E��V���H�9��0d��m�n���V�Lh3p;���7�����T�K�}�qp�1���鯾�ꅺ"jg�RpՓ	q�z����9�$K?�uf#U$ԿBB��6�)C�*��B�M?�<)0�Y��
hE�MnA��i�e:�'����=��Wc�ɷ8�j�t��������J?��s��z	C��0p��I�g���:#�I�i��?�:����!R�_��cfUWY��U�|N�`��њ��;v�m�M��;��\5?�F���l���Ѱ'�������VU{���Ҫ�V+b<��I?��:���S�<A��6�#%��Tn���c���U��lBT0���W��Աc��IR�z#�}�?�_:݋������O���:a�;����<���}>��+7E���xKYR߿2�|�k�X"Ӟ03~Ɏ)~�ӣ��r9�n~��>�3��t�?��B*��~��F�*�y��M>� <G���{W��[�g�k)����5�A�D|�&��c��R�����_w	unkVק�Ɵ���L�>�ܺ��)�c�k^����4�t���n���!�0��|/@��ٚIش�z�n���ƺKv��l����]81q�����p�+���C߇>E�$��q�I�mU%�E"@�l"Q�"�AQ��q�sa����&1��]�g;)�h\T'���D焹�>�&C0��x�<��(�Է�RD�f��5�a>�����1'�#���_(l=�@xe��?��}���kN20ĎpVo���M�q�D�%�o��	)!�7�T[�ŕ٩b�a�~N�/74&�W���e9�D���3�q=�o�7IU�.���%7a�v"5���_���[s�]O���-�nL;���s���Ᏼ��Y��}c�*��!��6~��"�.��3!m"�#�=��GO<�7��^IF6��K~�k�G�#�+/����E(ǅ.�6��ށ"lj�U�(�˚OR[{!'T&��of��c�j.]�ߝ��N3�/��*C����������p&�#_�ǆw�<�P��J�i�I���y�����c̯�3۠R���x���C�
ׇ��7no2�ݎU�3�]
*��H�nt�r���o�P^4�㊋5:>�Sf]�f�<�I1Y�"��Pg�+�<.�)�gxh�ߝ���viq��,�_=�Mה�x�{,).���>��G$�XqLi�zz��!x;����}���=�~ɶ�몲�6�_x��\A@��Ș/3�;,7�N�M;{��&Hg�����}�:
v�v��Z{�T��	�R�`���$�BR�L��'����.ؗH1�/Ӽ��w���G:��s�(�O��ǈ���4�G_��F�����WzN�-����_e)3W/2YAm{�ͽ���>�ʜPOɄL�ۼ�T�ϟ(�)�'e�%���W�N��t2��b��=+ ��w�ڿz�9Tk���W�ʑ�5/W4z�6�if�ꈔ����)L{#����d��ǋ�G2t^��s�^5;3��3�ܷӆ�n�|�����C0��c��A���p߿���Yfy�k�}�q�{�x����`&�xu�m$��/��}��G��J����]-o}B�
��6ġ�`rv��ޫyixO���B�)�H$t� ����azr����&_g��ǌ��)-(�Prgn��Ɉ�`T@)��Se D�킰_������=�׍��=u�.���8l�������4�YV�L'8U5I�'�j)c�7�+��-ې_�s�H7�a���{_8
�Z	9�=N2�����Kv��=�E�5�7�
�W����R��*�á\��0ZU���L~]�'���Yk�����\;-1��k,���<�n芰��b8J%ln�&�f��u�x1�!^Go�8�':�s`����@�AX���~�]m>��~�c��p�V9�0kؠ���{w�8���gg�d��g���]�-���S��ڛ6�g��%`u� U��nk
S�����s:����+�,Y���n��际��{y���[�y��ۉ�]��~��Ŏ���w4����ʋv�E�]]�&]��'�5��b[~��Y�����;=�*�	R8����u��֤f/5����ʖ�Q�}u|�EPG��G'���Ǡ݅�ؼ���ܰ��@M����#�/+7�� |�&Su~c�����t��e���v6�A��P�v����y۲��bCf9�'�o7�ϖ�o�*����Ƈޱ�_���)mk�9�D�ς��Sn�@�+]O�g~|��1<��p�KZI�����r�o��`'�a�Y�7�箸�íz \����N�Y�z .����a������4b ܆xO9o�����hi/`����轓Cu&g`�|�B�=�i��,N��7}��܋��;C��y3��A�7Lo�3�����f��\F�.���͙�0��׺��;�Î�ghr\g���2DVu�|ݺ�����ro��*���qI�G����qA$tG����Q�a�E��*�J��q����$t�^�scO���Ư���bu�v�A Gh���)@�8�B�i�\Sҝ�h㥮�3w!�*Zw 5E9�������Z�U?�OPp��]�u���wg���,��,P�p*�f��g��M^��H�"���4���@����f�B\(i2H~�jgn}To����[�ym�-pe�Ҍ�G�DA�[�μ��������q�޷�@Ǐ��*"|ޗ8 i� 	&�&�ʹU>-c�~E���YX��dXY�}��[�{��{<�p� �p��Q��j��a��Y4|#|捁nT��Db=������Y ���ZpM��P r�����#����E�渳�M��S̭i�nk�Ą��;C�S���|�nNC��"ZČh쑇�_�UJ�{�&�c�b��5t<����xɖl�/+N����gW�s9(�U�Ͱ|ew�@�.�N��:�k�w��0�\�Eoړ���?��;�J���Q>Y���w,��U�D�Ĳ��
�~�v��{���o�y!��ٕ�$��m�j�	ے5e���^T7��6ԅ���Q_��i����lh�K�'ޞ<� ���/ȉI��#�2dek�G: z���_n�P��J�rX�/�'��W�'y�o�!��CR����BQ�-��Y�����V~3{��ۆ)�� 	4���P�Uī���f{����B���-���+�S���:}.��O���?��%�9��+vF�����$�	���Sh�-��(ʪ�TKY��PK   �I�X�{9� �, /   images/c24ad21a-d149-4590-811d-5086112a7898.pngd|	<����[�����d�TdM����EvBY"��3�#JHe˞Bd߅�dϾD���w����9��>�)�}��^�����y��ʊ����9x�*��/@��'��３�����_����<�0���\ղG�J�ﮪ{�j��Q�+7Ԭ�:8߱3F�����Y��ޱ1泶3�$�1#�q��_�.Q�����V<ٖ/6y�c�O�{���v��!z���o姃�Cӯ�
��g�\T�:3o�L][z�U(��U;A(���lz[D�Bz׵[7T����V��`�_z{�{lb?�g�.nڎm�@q{����&̤i-fP�����n��|al�~#t�xi�?�|�.�\�ϊ��;���zE��'7]3]ݜ��C6Q�9 o����������H*�뼑�;߷dFj��2�)]���w)�������Pc�9a�%�� 1qMj��Ɇ�&�j%��U+����4Ι)[=�GZ�\[�W�<�ְ�?�c仵��Ӱ�v��k��]��S���.{�ZQAa+���:�Q��ʕJ�c?z�i�旭�ǕJ�{G�`Y�q7�"X5>92i[��'PѲn*Ko���3��{�b��B��" y��������e��g��T�����1}���D����)FU�x�<]��r<Iv^���4x_�?�?�N�}{s�t��O'�;��E%]f�2���u�Z�����Z�x��^���C��۟�NJMG�^��4�T�n���b�R�{��ӍwH\!r�n?�D��ku�׵���b���'���9���}�ğ��-�c_�\'�[Z�[��U�a ]��{�?�Oy�+���?�c��鶫ܚ�^e`�e�޿��ew����cI�T߿�긶d�r��i�}4�^��\|,�)O�.Myh3��jӤ��I*�s����K�$OR�U&Kl�����~$#���\e!j�����5����W�����T+�A�z̘��_+���֕q7Ԙ-�ի����
ĉ7mb�����I��b��]�����D�,��/�)�;��<�97�8����{��2Iړ��D*���Y�����F�ңƬ*���J¢�C1ckxL�̿�H�4D6��T��=5�a�b#��������N�*����D׫H�yq���w%�gc*E�pw$�vu�{ĝt��^U.zj���UUU�pҫB9y�}()aYXX�**z�Ei�B�FZp���vXlF�9��nT�KS�l���깩Hd�n��wҵ�:��[��I�^�n0�R����~�	�P��A���$�������ֻ���@
2TU����ZX�ԏ�M^@�g퓓f�S�Ǐp��C$[3�I�{s�W�+��/����l�,&vvv�3aG��ƻ��
����.Mv��)�h�����P�kv�ݫU������v�s�;�8��gCj���ix�w����?s持��9G1}|��ѱ�� �����*X��컌�O`���G�U>|B@����\�ԃ�4f�������^����O�j,|���␐��7o^�@H����51	���3�M��ܩ\�� �������ͯ�ݼ�y��'�/<<��:��_w[6���5�h���F�D�����o�e�ry�뼟�A 毸Ð�+h&�\]/:�C�ݖ�&� �<�����YCCQ��9TVZ(�qL��b��H4\ڜ1~�E'ՠ[�&� 3����5����}�9�44������	�;pV����šؽ������r�1N}���4_;@em�d��N ���n͌��u7�	I��j������C
;@6�L�Y@T4���Z
8�z��q!AA��+R:��.�w��Nv�eeg?G��_[[{�9�b(����$�r ���q�����~��u �FQ�b�&�������8�H��|*�(}?J6	�R� �Χ_�.n����#4#RJ�7o���@Jω�2vf��c(���Ə��O;IP��ƶLO[�+6��������Gh@�t 1��%�[Eg!�W�B�|� C��{^"�����p_0��/��B��<����4�w�,�㬬�H��A{W�ohvE�9:
�q��{52;G�
�SѻO9�����'�Ūՙ�+��o��ق*]0)4,l�V��i�,�}'!`�+�-S!��@hzffm{��$S���^uV���q/�#]��:ɨ���>�����ni`�+K�組?A��L����"j&C?���T}�53;��(�$ʇ�֢w���ţѻKҠ����ˁs�b��Vj��H3/$pd�S?�w�������E�E����wu���3Fح�T�qj#�p�|�u.�S�F=�P;�з�1��43n]#�q������Mdl��ðnvQsf�v��ʲң���i�>^�3�$Ｘ8�l{[�����[�������P�s�i�\����M��(;*$��q�3~��}W�N#����e�㕯Oy��0�H�I�1�=p�zhh(0U=6����P���f0D��U�iddW$���-�5�J'9�b�J���{g��grã���$C�b''H��s]�\�����"�9g3�"���������"���G��āW�,� D&��8��
�|-��D�1�J!'�C���)))�/{�U��vV��b�G�
O���H[�ڟ?��OEu���4�=o@4��	��C�x���Q48v��\)ѓj[;�+fm#Z��F�h�g�y>�ֲ7��۬��'z�i}{��9~� </��'2��^�t��%�5���q�Y]�$-��3;�o�Օ���Gw��u�:��?�k�8����l(���W�w�������TbRl��%��W�,��x{{����AYF��+;e�3��S�D�{d]p��V`KKKxl������H[Ѐ7o�zzٗ�(��"���&�(��{��,�ކ���\��*v��~�:�,�i6������;�P\^>X����Ԕ���R(������Ƨ	ESLLL�ݨaV�ȶP1;E�s����n�O�a�wa��~͈ :�L���G�41�w?$�r�5@gnm%3N���Y(�P��.3!��_�ྼ�2V55�����Xj�޹~�S�����<�ի'�liʜի�.Ah�4Sk��tuݼU�q0���HzΓ���Zx_>�4�9��	��5[;���7��� �ْ�������k߫��3��X�ٸ}��FhIQ�x	h��ܵ���{���WV�A��Pn����S���B4�heД�A�����ma%�_��X��z�ڕ��n�~�Js�|��ō U�}�����I���q@�@Ġ�$�>�+��B���H�cb� �{zz20�_n�z���ڇ��$^w-ZP {���$(���A>/8n��F������0�G8X��R�����uY^�s$��+gcp&���4����,v�_t�Q:�^�r��d377o��d��t���B�%�I����٢��J KW�Z9�)�O�D�\)6�����ITle���R ͬ���I�ėTm�������{k?Qq�_�.ۺ<7��9<���i�W����>5���)���k��W��Qn�^��L���`~čB�%��2w�`R�L�����9�t�.y�"��ר��!W�n�<����#�	����Ye�u	����͙���t���i���{��)���p�cP�f��^��0m=�@�AQ8/�L9��A}���ǵAɂ�yS�)Q����2K���UD�8��z �E���,|��cslY��&���s)�沬���J�Jr���0A!��)nh���/��-��&h��Z0H�?�C�m5�?{}�i0 ��D���FZ!r��3&Dܾd=B��':K�?䖵�vM��j���dA��{MW�Y�����>+�2)u@�.��O:��+\�_���g.��bF�yxd��LB�8�\������~,�,��Ğ���>��>+�n���Yе\cds��E�BJ:��==�:V;b]��Fq�LC��X$�X������k���I��>p�P��q�|������L����a$�2�`<Ey���ÇΝ{FV�gC���>g6��ϭB�+h��
��|�u���k�����_F�7kdG*L�:�	ܵAb�C5D����f��� ��J��O�����0�U���� �a\!hb �^��O����`c�*l�dՔj��B���?�8|+�cz� ���[g�!Tq 4��έ����/V�YK@"J���T2�S��5w
�/��"u��b!�^��˄�c07��BK�JYQ�$(�� *?���c�C���khMfF`�Kly'Z�Q���*�gX��"�� �"�i�[���!8q���m��,G�A����Tm��]6�g
.3� '��@9!'��SSS��|^䀍n����k��T@�չBnji]Ì�z�0��Z0� �{@���q��*���|Fs�kv��f+����G��.��18:��Ӊ�z�ݶ�)�K�!kJ��W(�Pctl+��-))� V�.�c����JP#˫ʜ��L>�JW�wXY��u�չ"PD�```@�'�R������J��%	Vϐo�9�!���?�]<�]o����A������D)��j�K�@㺣닏��?�ψ�A��RQ�cz�h@Roh�Ɂ./�����
̅
2`.��h�d�d}�����m;c�uqw���R*Ui�uYjm��0j_�B��gu�J��+d���OI�k]��˗jPO�>�.��x�:���.�(���Vd���.���9�߿���z깻44$mTS��ѻ/O?��ʂ*�i�;���`#�0{{A�(�5Z�~V�����y0u���x��3�#BWR�G�w'2���i@�i�,޽�!1�@����T���\__W�ݍ�3�Bc1�*A���;[��$�/u/�/�_?P&![_��ո�\���v�pS�֕
3����bB�����R_��������K�� }�P�q��bK���T �k���dH)ʠ��P�u�����=Hs^��5d�r�w������y4���Io`a�s��$��")��i��h����D�l�vJ,'���8VLh���	��&���.Vܓ�9��f��s���cC4!��<�x�J���@�NLL���D� �n��?Af\\Vy�"����LO.*)�pMń�`v�u��d���2&'�9��.��4>�#�ڼhj�Pچ�;��$
[�I	���$}�ܢy/�gL��{�M�����cj�u�<�Z��:��2ܩm�K�ͧ����%�Yl|����*<�M1�p��z�"h�hc�Te�CAT}��/�%�f���X�1|���%��0�y0i� �(���9&ff;�?��k��Q��ZV����1�8b�@��d�6�����S��/�s�n���%ƕ�P*�h���� ed�@�[��+p[2CK&NP�!r5>�Hܔ��ZDh1@vqۗ4�x|��|�
W��,*�ƙ@��J%M��9B5������V8�%�~��F�8�3'v�aXG�4ꞎ�밍����v+��l�AO��̦Z(�vۡ<#��t�bf���^c*Z֒CtQG�>�(�s鸟1�jٯb��À6�G���r�$�g��)��-`�Oo���5.��:�CA/̧d�,�f�_�-?�)2�22n���E�����-l�i?�2��ܨS�R�ዾ��ۜ^[�1~�'�0��h�S20�:�Hߕ���ebf6��664s�Ʒ���������'�h��"���sݙdn;�6�,�c�K|��C�U�n��u�r)i|W�Ŷ�.^��9����e2�8�. ��Hڌ�&�����RT�uf�
P��n<��sByBE�":ע�fg�}s0�7yk��U�;9p>�+��"iQ�_�����q�3���A��+KIi#��`���/�\��z�ﰶ�a�; ��,w|j�~��~ /�6��8�h���s��v���HV�dů��ϕ{��$L����Z���PVVvle�~t�_uRj�E;���ҧ�~����D�����kOr�8u��=&Fh?en%X_	���M��y6�
�@1t��s������[��v /Np���i�u %����l�uOcA��9:�pO��(�|������w��$V=:A��=&�%�{|\f6&9y�@�XZ����@���g�p�,7u���Ub[n�@36����I����؈���J���RbY�!Q��L����Ԅ����{���<�ϩ�����-�[�nK�D��Q>�\!�H����u���i�I�ˬ��C_A��Vz/Ǉ�H���ŉ���9W���|���HyP�R@��S#z���Ǐ+��^�K��)#�|MH��s�������Ό�3��=6W>����.��b���n�Ug5h�F�3PSQ!���a�)��2C��/@[4�H�~zj���P�ʜ}.��bA��)A5�@5\a�@��~�?U> j����}�����'�n�k�\������M��u��FJ©v���`X�[���� k5/�������IZ��\ � }n��3LoF�$��ϗ�7� ���yէ|��p��|h�lA/��vOp.Z"�C����ud�~�HO�\[��
�_�kLtf�F��A�p��x�,��н@K�������M���Eݩ�M���_#VJ�w�$��ξ�-�\���<�ovy�C;�Y�E"6�lw�~���~n����lC�lNS���HZL
��p|p�G^�l���"覐@�c�i�N�g!#�S;�ЉxG������7&գJ�°r�6�����X�����j�����6qms�����sk��{�Ԁ@c�����G��S<)b�����w�Шrtt���5�������Yv�����p�w���F�	G���m?��R1�b�	��^;�	����r�%�y�q1.Ï���w�%>�����p��u�Po>n��L�a#�Ǘ�����P���;B�Ϡ�iK�8���_�_Z�@�dE�7�l�yY����XUcE��XV�O��L#����W�L+��p�xZ�Z:;�_�h�3@ᕤ�4M#��C��1�o�;g�=0%��zn��{\@��K>��)�"A	����3����x߷=yP,^u���G�����>S����λ�$Y�Mk������g��h�=�U)b�8=�<�ud����s?S���|t�=3jw1�c2����E�h���X���%�E7,��$JҎ������/��PH��=���{�H��	Ǘ�mM��_g��<�E�� ��y�'D'�z��e�EvBCTY+�#�A��RTk��Ġ╃o�Җh'a�0�5a���
�{n���t'� ѧ�\��Mfv�O��e�y�˗�5_��0�Z.0<�l�Z3��7'>�q71�1:9D2�+���T6���]���J�eښ���;@�|vyCf$YrymD��5b���ё��Y���<�� p������o��H�s�v\~^�.dh�����Ab��3Bds?s�����{�,q̲ˋɁ����C5%�Ƕ+B9.K��7�>z��f$ѕ�6%�>ꖩaͥ^s��2�fDe��aAgX��K�b�?�$uL�&y�X�ծO��$Z�"R� p��;uw&�Y������,�M/�z����������Il�;`K5p?��b	@�u@"�p�d��	_��>WC�}W�q[�S�E�����=�ZJ�l�gM��H�X�S����؏���4HEd@PP� �ļ�����U�N{Y]��Z4zy��ƪ�Je�US�Mx=�Ի��"����!�O h��WX�O�J����:�絨<�d9�=rX�&/@1������?�u��r�$���xK�Nl"c�Vo���h�s�+I�j�T��G�
��F�~���Z��r�a����� ND*g;,���x6Ϲ�������F.Ӳ]�$X�;_�ĸ�f��4@Gd�c?��J����6z�;�T�<�!�f�Ag�G��ȸq����������@\#gAۇԎeR��$��)��,�0�i����CT$ַ}�:$�u���Pc�&����o�������Q�<f��#?&E�&d�=���ȣ��C�<D�$�I�)])OaG,e*�c^��B�jȫ�(z8U�g�`vt��%6�Yh`��곊ژs��܊�����N����(S#����iWb6�)�q��W�]?߸��:�LN ��6�3&���\]�\����kay�Tu���P�wh���@�����)*���~�*
��.d�9-� c��:K�↨���:_��l/Z�SˏFd��^O��C��f|ns�)�/_8�	Dr� C���M��L�Q���G̀[ﰹ���G����<2�~�qy��7�*�h�Szs�@���KtZ@/ݏN�����R��<��N���?�woO��Ѳ� ٙ�&,F����~Ĥt�a��P���TQ���'4)Va�Z���r�d��\��t�I
���V ��x�}v�K' d�w��D��y#��ߓ��X�=�Hi���]��a�O�la��W-^�:�~.��e�4���M\��;���H�@\��|��54��sG��7#�ݎ�:]@}��Yc�^,ɸ�,-�����l$N�<�E�V����\4���dv�j��#�����XK��:ǩ�f���tQ�g�]��e�-w��͉>/���`�YPe1���kL$�Ls�l���j��h����6gUeY[�5�&D�l�z=��q��2֪��ڶ̤p(�j��3�cb��l␼3Z�퀝���Z-M2ڜ�{̦�:M}����T���@Gי��d�������hֶ��+��dWΡ�9��?|8��T�4d���7]��$�DT������f�+=�%i�m�k.W�7٫��B���������5m�4n�]߻D�?6jŇ_P���o����gH�UyT�f%]釫�&G��G��2S�
r��:+�;gN�T��+ŋFZ΋�V�*./����:1�����[�W�+%饹�D�"�]�e��������dM�4�f��Z7�'=�y�ڽ?^�^�9��Q��c��nv�~�X����e�/�xr���i�b����6���hO�61��Y�	�w<<@�M0��ҹ��i'7c�=�Ī:q�뇈�ҡ�2��}T���8�HjB�vzڶ��N���T�xK�d�<Q�i�vٞI1�.����ݘ�4��c��s65w7�b���c����J��y^�x��5�_�~�h����k�@L��ai����m����m>9j�ه�!�9�rl��ˁ�K�g^dཱི�9E���{�ӊ�-�D=�ާ;����j,P�~8��N���	"��=�F�c�/�#R�u�<���b�OO�Zk<S ��ի-�p�kۼ@��p5�Q	$�)^6�Ua' �1�^�������Y��D�-��j"��Ŕ+~6^@�$�JE}��BOR@0�@��ɩ��\~�KBY�m��'D�m��m|i`hV���������"]YT;o��i�{�:���Y�g\����梗r�(K(�k�����R������r|2��ix~�(�%�FBa��7!a�F��ů�����ˋ�_����n.k!�y0�}�D��PY�b׭��іs5��3���QpE���k�H��`Z17r��{4�F}�>�6ȳLT=�s��2#'��
���T=�.���b����=ʈ����@���1�N��erP��;_k���` W/��9�;�"��d�������]hŖ���]}_�ş��M�&���W���S�	����,�t�m��)��g������cܧ�Cd͌��
��S�ɦ�.����2
2"Y�ܜ���
�Ǖk<�UZ\/��W4Z{��J�>:Y񩦻�C�G�|i0�xQd����r���qYn�H�zxuA���`C�'_�)����(���4��b%ވn�=p��a�4���s#A�� 4�KM�".r���Sa�}�7��oH���yes�Z�KU�vW����5N�\��gnԭ��l0��a��������R<z���>�g�cM�&8�US�''��4o>�i���4��1�?n�|���� *h]�R�_gj_ð�n�fw�Zx�O�������j�A�b�Ť$��^2&N||�C�^��x������<�~�����]��^;Y#m19�?~u�k������①��~���'����G��}*�n���%-������PUU5���ɅN�L����c��O�cܸb�&SV��$�7z:����̢p�>��sS;̌��:	�ӓ0�k�ܨ1�Nъ9�$��?�V\v��̀�O�|ov��2�5�ڕ��s�J.������c�!�Ӷd�Z���F>�sl̙��tO�k�oO��$'��|nI����[�e��.��c�[A�����b$g�fb��S�2��>���X�fl`K���c��J�f�|���3v���d��������&��N��|��1�3g^��K�p�zV��ս�b��nx�='@f� `���`�=F�?�9܉���|ȋ����cB^�	����*�%���(%��ٝ����/��b�!y�q�p[Y��9'�'5��u�
�
@�����B,����ş��,����]���͓z��dfx\�-]�@�I�	O?X�H�4��L����6\8-���s�kLmi��6Yb)EWr��V��|������g��E���;�3��O~�]��ED������J��G�${�5o�ʕ&��s���mSЊ���=��n@�@����\,)&��~y�>�����0`��9�-3��߅p6c��C۟���Kl�%�%+F?����O1��M���;F�_�M.��@?�xuw�Iu`�����=���C_s=+����h�8c�b���tQu����!�#"!�����_��x��gwT5�M�.8��Ę��������o�����8��I��.�-:��ڑ�4̾���p��R��F���4��Y���(�6$3:�8��S4�]��ɷ<�"�8{u-��V���=����Z��w�9~�ҙ<]M-�=�����������Ӽ�/y"9]��C����7P!�o�	��Wg}�ɾ$�,��HJ��	�~���,�b(�e��'���Ư񋹞�Q���`)G�,�C߂XP�Fa��Fr3~2ًk�޽���:P�(�/�"�:ۄ*4�?Ħ1?jxK����װ�zX�Hƽ> �;i�V��B]�uYFϊD�������nd��*�t�]V��T����ܞ��G��b1�z��!�D����3ړ��ϟ?���G�s�i���l�.���YMb��!�g��FW��upI��H~sn'W:ߠ��`�F`��=�������+�r��8#-�2�ʭ��~��6�꿖��Z��ۻ�^���>^�ޑ�~���c��s�r���>Q��/(�Z;��7;z%l�yC�J��=�[wn|Kv�"&fuU�v�*�c>r�U�nZ8�"r��X����.Dn����\SS���'k�$V
1����rIV��﫟D˲�?*NMM�g�d /���6�Ɗ���w��]<<�_vC�T��p��.�1o�G&c��/"ϭd#�$�������O�M�����^��"""��^S��+^���tt�S_`.];]&�r��E�m}�����UJ�/Q�ur3P����4<p���xJJ�<��F��d�����R���'k�R��Zap�x.���s*A��O:�����1W`gT�i���h
6z��'��.bF��c���xQ�����[�I�G��6�|�1>n��<������B���Fdط���d�����cb�{��D��n�d�`w�-&5\�!����CJ�<(e,�nL���n����%2�����Β�@+���c�k��zg9�>i�spɑ�_�� ikp0�PFZls�
�ǐs)W�?�I��K@��izX��>3w�Ѻ��v�Z�܂�Y25م�)EEIi��b-�|����pv}Tl6���k�vX�R ��!r�A��:,�%L���p�b\w�J)��ݽ����m��=�ߊx�:��(�T�{.u�~����[�ek+P���9S���1$>�4���@.�c�a�t(�٤��w����`9��$^a/���i����+�P��eKgX���P%)�w0p��I�e� �,(�d�i.���v��7ׯ��|ܓ��$z\���h�)c���f?��R�R�5�1F���``��%���l#���a�QC�����7�)N�es�/��J�{�w��)��������"IzWȌD�m��oQI֭_�\o	b��[H)-��������z�EU�q��#�md� �'X����^��E	5�%u�*$�K�������?@8M�����,Z��X��,��I�����l��s>���p��b����?33��ڝ�|�����G'���eH-�������3�����lM!Jg�(qw��/����X�ŷ�G�X,���P�5�[T�S��2���Zb��
���XMu a.'�܃k��sY����C�2-����l�?�>����]ԟ��R��k�-����\�)w������ܮ���1毎��.v�Q>���+IIgd�E�zU�V���hd3i����ԏ��۟�5�_?�tKsfeb��J�k1w���?NW%�TPB �MMm������bq��#W�&K0�5C��1Dg��<��벿�F����D_s�=w4����s���h޻iV�#�>o;zɉo����ڏ�yj���W�>7^��>���J]��N����g����o����6�}d��/oR�+�r����ic8ܷ�(����U.�9���;��WSsE����,Ī+��F#�J��MM��쬩^0��eH��g3�����[��,8
���-(+�;--�h����%/��}��Da$�fh:�{�	�.�l$��g�z�ǈ�ħ��
Q%$����骼��g��]���>�ȴN8�5)�:�j�65�nzdW����,�{n1X���V��Ӟ�;��XiV�Zn�;�����x��WX�����	�`��+�59.���895%���S^�N�X������lkOBs�Ww�����˚�Hw�j�[��>;�M���pk]{ �cnv�~g�';�Z��0���1ړ��B��*P�Uv�!>l�qw���*1!��r��y���wG������M��_�d�&k_�շ��>72��劃\x&NMмv�P�˕�DSSS�L]����R̎5uSs㉵ð�����.���>c���.�?�ѧ�nDqll��R$ւ)�3�T���\x70�GNj���{�b��Hr\�b��}�Rj9�����`�����&�v����S22��}z��L��
5��xP@|A��M}&�R-fVLn8G��Z;�����}�J}Wbv���K�ƍBɂ"ٌ'��QXN�#!V�j��6���]��._f�:�2���U��?��q�(�����2��sq8K(��K��Z}���"�':��f��7��R�4�P�¨lSN}���2q�ɇ��;�<����[η��'7I:6�x���i&����`2>��p/-����0݁���9�����Q76623�~�Y��W�?_�a��N|�%��h���:.��h6[�Y���-�0z�x�����4������'�ً��n2K���?��h!/<���7����j�)'����W/d�P:������d��Ds���X�2{�����dkGN.Inmp���M�2�����A���5h�C���[�ŋ��!o�`&t{eaa����
�=9>~�w��5D��,v0��Y�c�r�v>?^�Qxq-�H��u��!����}�P%�o ��r������C;3t�YX�~�fS���yrA���N�0�Z��d�W������,Ԅ����]q�Tl��N�a��uX�,S��� �TeN#t(��%������Y��<���}YCk�����|k�F?�[���ѦR�<���K�^���ba��]�2J���t >�~0�"V�2�THބ�?�����Ik�K�G���s{uR'iu0%?�������ġ�{�������`ܱ�a:0,˪��9z	L�����ʷ����e�W��V�vHSJ�)��w���Է����vuk��V�1p"��{@�D��y'�{vc=V�[�.i��������ϭHQk�ߨ��!X��g�&Ds�}+5���<և����}x�7�\ ��q���{����[!����.���̼�(+�_�2���D���0�w`������B�%����ivbE���klP�df�������y��w��YtL���qY���/8П/�ok�w:w���ܾ�;�LZ�H/v�^�ů9�o��ԅԧ�l�������/�_l�Y��M��M�=�۹��� ��e�0��������耵DW�8���;�QLP��L'gmH*�+"��S�y}R�����x_�ǒ��!�b�Տ�s���y٤������?D�����*�q	u��׆j&�L� �Oj�	ܕ�2EҔ��i��~[2s�χ�-��N�7>�QM�42��C��P���xG�R����W��Ϭ���2D����F��c�+p��qw��hh/OC�e���N�uH���:���;U�т`Ni�S��ߐ��f˥�x�O\��.#_̀�S��u�E��J�	�u����lf�]��b3uu�v8���Ӡ���D�K�z� �K~)��+v{+�����wO*�lO�޾t�W��I���r��K��B�%�D���k�b����M��^�X�d3DsU/S�7ߺ���[b}��s��J[[�<y%��_g�
����ish��m�1��A�����lS���)=<`�.�T
��2]���J)�$�ZދՏf˞)��c�d�f�X<D�s��������ˌ�T.��z�,���:���ƚ"���Վ�X[gZ�2 K���������#x�K��ŋ��!��͞^��¨�/���m��$w�JG���Myb�|�{��&�������Z����dw}c�cp0�0���xK�i:���l�J�[�S�6<w�Y�׏�S�--�K�mYb�XV2��s�skf�h�Y}�-`�x�M���=3��9l���?(D�1�����S^	*�>�p�Ќ.���S[��`��2����32�,,�'$$`ݗ�M�6�{��]K�˩�����F~%�H�S��@�[�e6��I6�M��6%|��EY������k��I���W��h}��]�l[V�v��^���+S�l�l�KI=|�zG�Ǐ�$3k'V�F�-{� �F*�zz{�T�DW�B6�_�u`�i�nzOOG*i[���7�v��4�K�x3�m����>9��SS��8f)Пo���dt�n�Ր����.5�Ί�EE؃�޾-��:�#D���>	��*�M�r˞7yy"�yy�))��� �����
p��v3�����	�x��� ��Ҡ$G[�ni�:)w��N4�cRaN�S�/z�o(WrF�Qy��Vna!'��{w���^�h�4qX���&]?u��eȻ�Vh��S�M�Ra�M��R�`��W~���}{�wWܝĚh�s���8�����QLDxK������� �HЀY�[2OZv*��:v)ɰ򯼐Z�<�v`�@ͧSn�J�����$@���,�w�����K�n�^�-qQٿ���[�����@
�8��2'���n4��#��36��
�~I(Y�U}Y�u���j?��5�I�1m?�h`$�G�%�}������s���.�B��5����W�ͬ�)w�<��#��&�����f�E\��okA5q�����~CV�V�<V197'�MHHw���f榽���g#�V~~�k�m�::�[ ��^j���m⸖����v$*��1R�����v�=�::�ŘK'��=q�k<��|����1!��7��7�ҹٺ��_t��M��i�p}��!��\�!�c���-�� �!�qnH3��]+t�AغUnǮ�ft�-��Xr�H���T�Lxd��:{C� ���׮�3ߧ�J�Q�� ��\�P��4��LQE�ҮN��(Ǜ�C�C\y���
����O߲��oU�����`e���<
DPJ��݂�+�o���K�����%�2���E���@h#�%��!/L2:�;��$��uR���,�=�C�R��s`w\���owo�nWuEK�����:��2��n�������7h��{I�����%Tw�Ck��S��~����=.�O9�n�{k*d����5V2������IIg:����s#"��ζ	(? 8u��Y`e����lT��OQ�J���p$��ި�Ђ�D��.uǝ���G�`���o��\|M�$�'�_?�7���>�)$!a��+�,/��6	{��a�5�G���?a`dDk����7���c�ofIl��~q�M�wĤ�>>(F��=�fW��ŕ���g/@���Ye(����s�|yU1V���j���������l��ߣ����ICPP�UD�
�z������^�~gEY���E=����[��L<J�0���Ѹ�����@����[o/wlS�I\5���"Ȕ�z�	}�\\n�|������/�b��^��D��h�r�n�Y7�>p���mJ&��>�]�W��Y� .� Tý��lkI�]��߼���@�������(��Q=D8�o����9`�Wv��D�lX���L%=~*�@!��/?�`r=;�o9��t���D�b����m�~#�6k��B8P؃�����bn�*�Jr~]���Ia�����?��#���ڑ�5?����eU=�$���Ϻ'pA�y<�_��;.X�����Q�(���|��|}n�A3jx�I�H�m�D/_d��
���8�t��*7�<�X��9��S����@^�U=���9�,j�s�?��h����w>�����;��|�����p@ֆ�R9��}S������/�
��6��yWܴ���/T*��p�$]� �����q:CM1q畱�릾~��BD�[�4�����:yQ:�� ��uV�d�=Ŀ溬��Ő��+�}'����eVaȿ�,��a�$�)���O��~\�W *x�Y���\k\�;�Ս-D������2�>J��y�'ҽ߷�m2%���^��GfT�&������>%ٔ��VU�æ�z�n��
��g��s�JIK�D`ʪe}��p���"\!���sk\�"�Ce4�UIoq��M��xR?G�~р���L�4�b���t�\M���b� HΩ8r=����rtvn Be�̽z���F毝Ck��3��i�Ž~�s[ڋrE|8�z�,P����_�����@F(��%����{�vS_���VG�H!\0��c�a�^9�1-���~���JO�YpJf��������L��/�j���#~�'{
����gm5 ��(�K�͊G����٧�;��b�:ϋ���uu-�25�`���t�<�&V��ߍ)n�!���U����X6�'����6�U���@�,�������� ��'�9�N���&���{ڨ�~N��W��5�|+aL�������Z�x�=Hw��7�QWn� {i^�(�`��WF�{OM��\!L�׻D�z��4e'���;���c��<wA����h�?agH%ן�����b�u���ݽx�tLY����΋�s~��������LN��=�wz=C�|�k�<i�%��|���>�ߕ����_��Q����G�(?�Dk�e������ۼ<P�I	�����2���~�1z%����ʚ������\�;uh����g�^�JY�@H���i-��_#�3n�R��^2�əT�՝�Î&��ޠ��`fbRVS{q)��9���cc��?R�89Q��|�X�Ɖ:����a�nwЈ>|����u�o�n��Ԝ����
�ND�zGGa�gc�0���
�r	������w�����ɷ���܉T:HC�
uR���A�	�J<޴�p�wI�~P� m�q�se�l��&/ߠ����uM�+�5Һ,�}+Ĳ���	���݈��C�5Ogı��٠"=�0����g�/����,�_G㜋�2�������;��3J�Mߦ2˭�e�s:^MM����)�/Y�$�+,�*_�\}uT��7���(J� �ݡ" ͡[I��D@�;$��n$ҝ�C�>���o�g�?�Z���<{�O�gόq}��;��Û6��<ܞ)<?E�wǲ����e<�����BE�5p���95�B������	SSS Ç��M�=U���������Wx��xа��
`J�䰎�[4 ) ����r?��P[��٭�ン��u?����ek�`��G�ϣ������k�wv~���%�ýh���E="7�2Sc�����S������ەU�~m��r܉#y =cx�O�fJbx��KN��՚���<�~9j��țD#�����aQIR2�𡡡���}�pB=��@V�{!������/,`��J�'�5p.�������B(hH[.��|�rKe������?���D���릱֠}�>�9B�m nC����s�pӉ0zI+��Yz?�jL��ZaႳӕ�v�sk@��o���A� ����p�O�����@f��X�7��E�or�x��H�9�
��/��b��M�u9'η�ܮ�0��b٬/��S�.\���<�	C��5��(�������*U��nG8E)Є�]+��L�ĢO���	�cn�VU� ��ql��f�@h4��i��"�]���U7g굼����"�����G|e{<���O&o~��X	�h��J1���}G�ni��������g�Da����������jL ��[����mmq�a�#��1�\�]̪{������b0�g}��vo,::��w�T�Շ�����g{]ADM�J��V����{D5:*�>a@!,�()+�BrG�[�_^�"������.o��^�%_�@�1C �(���M�980�*QJk�YI����tq�y�vl��XǴ�J�����Ȱ�eq1�%���hQ۷��)ƀ�I��'�B��܄)���^�ѻ��w3�z�n�H7i��>e 2�Qfp�_}��PA���/1J�a�ib��|(�f����N�JH\H�f!�rゾ�������f��w�4��a�R�4H�-�2�~��Cs�w��>�j�D_m�|���}�A\R�E��D��I#��d�A�?�<5�oF�q/�ɓ'�}8W�<{R�R���[��|Ρ���������d�r;n�m�j�i4{@/��]9�D��/Jw_�F<�-�Ȇ�v+�ރ�	K�[�,�\S�`զ�DD�\=d�w�5I���>�WS3����)S\(*�T�B�4���/i:��Y���uԈ74>n�-c��ء0�<��t��U1Ka@ܒ�� ������>ݡ���#�8^D�N�|��l�M���7ѿ���5u|-CBYaސ�Y��n�6�����b��
�֌\�0��vr����'��U��y&��d����MC�@\��>�����edd��l��n�fq�|gV5��O]���z��wun��#�쁾E���{���28ˡ�Ŭ����>H+�2�/�1e��	��F3Xᩳ[���]S/�l��B7,h��Oᔐ�&�����\����~��������s:��Ž���3<1a��*Y{������]A2�% �9-�tuuѧW*���5��l��	�4p#Q�����q��<\�n�2�)#]-8��II���3��]�r�`�#J����=����T����p���A�1Ц�:pf�tu����x�޲̀o;��ȳ�yK��f�\\ٺ��=׵�-�&D�M8�`sV�9���2���/�lT�ю]?�G*\�{@׹��=6|�I�=�#�;()�1	/�������5��s�sQ����O}J@@c��e��냉G�t"ޓ�ߣD��M����K�q�أ�	���ܷ��\I�
�Qܜ��	H�+3OAAy�__?3:=&�'�vV���(1����P�^h�\v999���Ύ�I�'��������]��j�EFb�f�{�T[}k�;��A��IR\�'OOO���hiWֵ.�������<�i��N]��՝���B�5H<uJ��fR��"�KH�>�%�0�O�\��ooca!=�C�5896���_mT��º:M��W�O������,6O��qm���{�� �=J�&{�-�t�i"s;;E��5%DfP�SXX����U�f#�2X�M4���¦-��o�,9���Tzhh荌J&r������NE�j�L�ĬuԅPc�7��(2�l����1�B.��+�O1���4���8�ͩjx����; w(.6xf��4��/7O�Y���UW��B��\�4--ME`y�HGUS�^0��_������u���]b8HN������=������^Y��V�?���A��Ҫۑ������x�Hw���3������"eyJ��VD:��m#���r=��fG��x�s+��@%�)r)��0A��mB$���&u^V�/3U���A�����Ӥ}¢���� Ozn�C!��җ#��t�z�ƅ3����Tf&���d�3�Q.�Y�ҷ{���U���L�AwH���Sg����X8��M122"T�%���\&�D�cVM�d��^��$)d��#��kU���l3a�~�V]+�/	�b-55�2���T5��N�[ ZC�AtE4#"�n!���N�,q���봵���s�ׇ<H�#��iH�r LO�7��i}vdI�S���^
bG�)��ڶ�k�ڨ�t����!�kZhvF�)(D�JJ3��ũ����8��V���
�6cJ0ގ�lZw����n<\�V�2��60(�P!��jm��O�3�]U�Z[[������ddD=�V�L�~/ј���4y��p�^���I��l�-ˊ�VlIs�Po_�UR���[1*�+'�ȽxR�AIL@�&!)����X����mF��a���JtmE��-��b�] x�GAM-�����S,�wۗ���������tA�ă��q�" URS�T=�lC=�w���Us�KKK�#()���l����TO�r����a'�y�wz��@��нcϝX���4R�~��������M��ں�a�O��3� (���Q�bhXV1p៩�πA�t�7&����w===� -zB7�k��r�R۸k?�sY��-�<�� [�Y��@�J _���Ǝ-�-8  �ALCC�q���1�3��9ъ��Cа�X�ڬ��=�0@gO�*ڴ�j/N��վIL��`c�Z�<Q���m�5"P��7����ܜ���?��͢'al�&\OE)sN��\<z�?��˶kC�4d�6���������ݒ�ڲ�e��Ң5�:J��S�nJ����c�}Ƀh�`u�[;G����˴��=G�����<9�w��s�wNa!C;Z"q�r��D]���Hc�'��ke>X r` ��ft���w$�5��c��:V�u���pj)(dЗ�����j�b���+t��,���f!����$��fm�*08�V��Qz�-xZ6�5��i],j��D�cP���$ۚ�C�p���Ͷ�V���E��bt����������CCZU�\Md�����8q��&�����[����uw�C�: ��U����
7مE�	
�$����R�d<��1�D)c�m[@2�'ݏ��3�>bl���jh�1:]	=#hsSAZ:���[�N�g�*�gi����6��^,�+ ���㩐WRʭ���	  ��.y׈�:�k�G���ʊ3�Ʒsk�R ??�
�O 5A�$z;���P��"P;C�����0
����Z5��5*O��I�'&l������ς��JLL\�������Z��v���t�����z�4������`E~H��Q�$�te[(��T���+&����!�yQ�`�Q Nudk�y�2�� v�@�t����IX� /�����ǟ%�
ۯ�PY����az}�,w������!�<E�8���[0�{�qڂ���4ttC4*��描�CsJH�i��((~>	��+���� ���\G��5�� �1pi"�Fvv#6�(hFF2B{�ee#6�" ��J��ϗ�h<ݝoc���f;OA
H������:�SP!�)B�*QUUUC��cc*��6��A�۫�T��j �J**V�ݮ�K��@��P��S��hk���=N[��?<���v�砄���cb���������o�* e\a��[(�TL\��FF�E�$>>>��������&3�@`�!��}I�5�B*��;%'�������?��<P&Dt���~�r�n´j�l���'�~�Qh���(b궶�e�3jf���,Fm<��j����g\˅ED��۫���i��ˢ�:�?�����x�[,:�V�Yht5s}l��%PXmk���+�y�����;ڝ/ؼ�"��$�|�.�Q/p���c6a�Wq�訲T�x� p�V�k�f��f�"A�cl�x����rs���TUQ�<� ��q�����>U.�d8�))|X�;6CEJJ*��U�,=p�������/���;KO��  ���CDIY4"=���J{(i&)j;LR2�pc,(��DW��2ӉLP8���kv���|�����?ڜ�U#��L�.3�`p`�:��qic+Ϭ�s�sX���SyW�Z�S�+�+ӻ!���8X����c��w�敒�ռ�3I��O�B��u<uP,���+ڽ�2tŊZZ�W�;�|??����{�x��ʴ�]��X*9�6b�G𷫕@�zM�yK}	�8�Xw���8�&%#;�}�����ʟ���w}��M0�a�c�uW�c�&��a�=��d��E<�x�%����&�@W�M�& &��N�,ۈީ����b��f%+*))I���HVU%&T��g^�Z)h��;�3up#H�n@ۚ7k`&��Fߺ�*��G�^�����r2�5�6�@��0PSG�G��$VP����0��ܮä�_�(�$��X-�C�*�1�� ��x�/��x;� �\gI> .TR�
$���2��B�sf�i^�ӈY5��9Ry����=���뫍�6[I����Ah?
��r��Ϸی���?B�F��+_����xs;��������P�/tI��r�w�`�q2�N��jG��3�O�PK�ݒ� ߮�O�J�d8�`%����/cu�9ĔN�q����k8Ei�������V�����l�6Ӵ�Mzf���F����r�`�=ю�j@A;{�d-������'�L�Hv�!��y�Z�)>�N�xw<j4W9T
g5��[Nr.x�=0��`s���	=D�<��J"�,H�P���󄑑��qM	��\V�M�H���u �i]s[p��IC������E�˕!����Ț�m�9��؄tA�ƹ�E7�M' �l���'.R�u>����]۬��}7�$p���Rp$udG�y�t2{�Uwj�Xyzp[L����J��7! mPVn�����h� �J�>~�+F?+�[��϶�4���8s����w���5�<[��T[@�s=�����VM�g#jz\�)�;q�
��M��>b��3�#�7/�ϕ����qo�9�70���)��c��?���Y�ag�X]_���S���U��)�Z��������I��S>��O�3u"������]*^��S�oӄ�P�/'�'�0,~�@Z���]�da��\���&�����m���ݲ�t�3�0��
 �`z����aU��ʜY�ӒZ�1��Q����5z���խ�R�%���� '-n��3&~bbb��q99����na b"">�OrA"�N׌�O{W�m�ˤO��Wʈ*�t�����n����a''��K�A�N1@� |�o����t��Qb����TUU¥��Or1�������߬� �ajjj���������@fF/T���g�������ߒ�F.�'��DM|RX��H&|�ޔY7 ��.Fн�l0��5�@��o�,��_>,3�N�h\-)B�X�wjW�]�N_?3����u;�x���L,]�R&���Z���ːz�?ȀB	���^�4!���@I�!"�� �C 1& W��?�p&�~�@��d���=Qč�[5�5ya�Alo���aG��:l�Y����EwB��|���hH��M�N4�v��}{��A�@����������S��*봈��F��e�V�Ȯ���5/$�y���Y�v���������*Q����}�$]�;Mr��ʈb��6�	�rPߌј[�N��IM3Ԉ�ݝ� '/�5��t���W�(!�r8b�\�L���p���۟�&�����"#=�E3`'�0zA5�QQ,�ŋ�"��YYD��h�����6�
�'�h�t����ft�������d�p=��?GΘ�X���¢����cEHf���#r֨fPL��؉�L�8-�ݻh��V�P߫�V�`��FKK�$����w�U,�f��ns���Y6��0���N���3��ҹ6��f�}e)+��g@��zV�4�S#33��r��yy���]��_�჻����0�u��oh("ԟ҅?�M�<J{`��|�M8����lY >�S�6C6�J6�s
���S�1����S�S�


��8�__]f��E#�- .��|x���8 X:�q	m�i�z��U%k�"(��sͣ���B�������Ay:�r�<�Ң���$����Qw��ͷJ�uwWؑ���;[E��hW9���n�ɢ,~��{�wt�>�[�ء>�C�S��o*DDD�,���i�ɣ(�Z��#/aC	8k4�4W��~����(-��k`$_������8�[u���W��$����(�%��*sM�(�K�\-�U_P��v�/B�#��/��6;7��_�E��o})�O���g��qʌ����*��ʷZ���`^�8蚧L����C��jq�]�nT�4CS�i�Jq[[f�px|jD���/K���d�*n��v.��Y�ۤ�O}�F�L*>�FI�c�%sQ��s{T�xRX4Y�#�FE%� �gh��C��Lk//N�k�9(
QQZ��>�qp�{XY�u��Q�YM�/�d�{����<��Vl�`���/xX�.�:T�?�A�����iCux{8fX�^>��;u02��A��Ǐ���šY���o##� p�7ųPh�����99�h7P��hޥ$�OCx?����Ggt������I��1ޠ�G�<�ɶ��>&HV0���L�� 6n����\ZFFF � 3sj]]ݍ��W��Ը�',��7>{���Ol7���c ��4�?]�EJ��iK���%�9oz�@���d,���"R1���/�N��1�6^��L�D*�<c��<�rpi�PU ��ԑb�u���g�G�����E���ZX���##F�ḘV�E��P<�)��8��ok�w��� /��//W�,��)��7������@{���g4l�
nK[Z҇F���(�Z��ׯP7R~�-%�a�5�-����]0@�_}|X�Ύ�*`��� r��ϻ#k��!�u�\Y�"XQ|�|#�o�b����'��w^t�2��ASFָ��@	�LZf� ����'̕X�و��|��
ј���O�o��R�ѹ���}5wQ�S =��z61�]Y���ln^�jF�)gm���q�� S��]����ܜy���6��;�G�^�G�s#�F���k�{y��k��<n%I���eI�e�9]�#N�SS�D<vO��c�Em����p҄y��M�q��!=�f%黫�IyP  ��.k�m�7?{���, O��`%�,��g72 2J�^����z���3��U���-6U���(�	H6V֧����� ���0�&�>��3Ts�����j#
�L�+�IWj��.�Xh��Ȓ��;�D��$T�l�˅�W���Q�!�*���ˍ��f�%(q��_ѹdD��VM��ep��;YU���[P��1hڸju�P��88��&�zhd��E,��R.n��yy#[��I���߿���� C	 ��6+!��ֹ ��;�i���f�rK�ٶߜ���n �q��A�%p�>�?9q����Ew�6a��s��+)E��wEgB' N�~�c�钠��>��`� -8����k�*|�N+ݫ �V\b����2�S��
�4 ��+�kiiͦ'GlZ�1�1�߹d�ކk�߫yb��V������� �K�=4x����,6'������ޛfTL�;q�y�6+)�8�P�"4HR���ۋO�\|���d���t���j��KAf�Ghh�)��\�5{�VKV)�����ef�	\�t��uӻ�m�|sWq�/��t��s�%�Yh�K���7Hr$/�e��y��O'
6>1ԟYI�9%<<1�n��=^��$��X��{XXOǐ��PM�rs���^B����������JC-�͉rc���u��CE��瓕�N���l��.M����e�	\iP� �П?!��Tʪ�`c�(����� �Y!Q
Ṁ_���\
Օ��^��UQv�TL��t�M�ۚ��ы��w����� /$�����ڎ�8	5[aI�I]6Y���[䓓���]�SߨkQQ�׶�9�ʳ��^5��~5&�yR�	�Hy9���<&;�������-,� ɮ�����m�Im��O���d����g.k���է�33��?�}�@�Q2[||�X��IsrX^�O*��bY����� K`8��8��M$[�Ujk���UT���4� ���HaG���Db������E�a����
��É��� ���z%g#󣢞��c���W3	��7J�Hɘ]~�$��2�IX����F�xȾ`���d����AoB?�y�G�T:�����gT?5�]\��w&����H���:�����$��UA�xC���TϜ贽O����욛�Л���Τ[,pl�Ⱥ�d�KV�͊��ܮ�l8d=9�vSi�y������������	�g1�<<��'������c9�/j4ݎ����/7�-ԕb�w���a��d]Q���d*�z�G���B�2R����R27HH�f����6�=$V&��a�KT��!�<q,D�,��m	��M��u���\W��"�>������	���Z��؂l������|����e��O>�\�p�D��Q���>��.§�vvXs��֭M���[�'�J	���pN-�����/qp����:=��gG����BB�T҆G���org��T����Q7�QsȠq�.,-Qg�}�MJj��u�=Y/���F�O2��;�_ll�nMєfv�����u��N�i�'�'|8*!��H��w+���Μ�R�����H��IH`��K'�R��2޿E�F���C1O�e���/���.����Ω/*��5E����[��Ta�>��'��?z���d�!���Q��?>�k�$}x�q����� 7���F`�����G��`�<��� D/F��g��Ǭ\��ȝj�^pj�xm8�^������p��Y�˗�0��L�ON��Ok>JRG����հԗ$�C7�jb�n~XI+������(;.m��C$r>RI3����Yy�*::�K׳���!��NS����/��ܺ��[n۬�}%�lب���O[&Ϸ����)B�A�_�m2���	;&�2�r�F�/�܉�>}46���,\����|��ի�{��k�/]xyx�
��J�>6�II���g3��˦����\�u�_c		���~+k7>���۝��+�kn6[�w|YX�5D ���A:����V����'k�3Tq`` ]����m����Ą�2bt�g6T��q ����3�����̷�g?^�e�2�t3�+p�%��:���ѧ�\���d?��E������aZ�9���p���a�J�������$��-�
B����{n��J�퇲�{aܺ�������)"-���������X��%���夜ǱcU˲(;::v����r��ocgG���w*-���f�!�F����ϩ����&�"�\��]�bX�t��X���R��*rSf�/�Rc��D.����P6ֻ�8cgO�wUKlIt�[xoX/���j�I3B_��g�Z�y}��=b�^K�}5H���N�m��Sdt�{�Ę���\��B�~��\�C�-�j�v��P2�����[՜�k߃��IH\e�^���j�l�ۂK��iZ�l�e*�[=��G��@�d�DG�(a8����� dm�b�9�M���뚱��	�\\�e#�XXHKg��䡬�KY�á��	h�,̈N�LB�H������@jzY�rjˤ�� {a�y�F��X�=}}����A��'W�+�����D��K�#�r�ς���gز�6�݇�%�{Թ'�=�G)�`)PW�N���3�����_0�|)@U�e-�R�/�̘����쐏`F+��,�F�%����#T3�r���լ�V9i>o�i��YR�o^4c�t�S�����Zt$4@g2��u�k��?M �!*F��]�h����8�ʆ�Xw㑼PE���,�`�Oգ'(������ׂh�;��S���t>��P���ss�?�����nc��������ϕ��=z&hfF/�-�� @#DRa��6�Ͻ7uwoo/bxd�6��&9F����O�11�������l�11OK5���72����W|�ƳDU(�U��K..�}�ς(���q����+���x���F���X9	9��4�8���S�D�٨Tl"����\/��U8��o�h:|��p���T#G�Zś)1�94i��-FfbG�[�|AHQ��Hu����g���5I������*׹86]@�K��0�-���������Q�*܄]g�����i����]5���J皽�e�+�T�̞}tb��^�"!��������wo123{nm���������ӻ�[��I���:�..5Ђ���)tfNM�d:T9�������3���F�"_�h����V�nR��V7+' ZI��*c6�ޠT5411䯡���gϞH�^�I�;��c��}�B��Gs�A�N�w5�)?�đ@0���(aT��D
fh��}���1�EJ��	`�o�߳MT��
+���y�mE:m!aa�X�Zu�?�i��^��ވb�*ȫ#��e�Sfmm������p��
*�?��' �V�P�a��ũUOR��ݯ��}]FY�W��X+�777�j��ºۨ���1C��"Q�S[�߿�88(����KHH��:$GD�>B�����7�w׀��ٹ: <���4���d�h$�'��F�-(b�,r�w��5��o�g���f�]��Ҩ�i��̈́^�v1ͺ=�,��Ofؘ'���"�)�;����66�iii2������}#���FV�U�������a����Suϣ�����P���/�I�V���&`%�\W�Y�Y�����蹊��9
�;��� _	� d��'���J4sKUz�6/�H$<TJ����,���Tk[[�$�g�L�.��z[A��~%0�:���r.��ޞ�x�2�vp���q����[������Z+����8�����퉾� �7����T@v}d��g/'?$)vU=�L@�{J@p�bk�Y}���
�!z��.��-��6��?�ý����mK���K��K���cʖ����`���)�%�dJR�Xbo��d��o�����;m�'�n�ҹfo�]��K�X��=!��T�v������]����?�b��������`n|r4/*..W�}Z��=���	�6�󵲥��v���h׸lٸN���Ց���$%q�N´!�a0��w�/��5��S�\Q��~�	j��+��?F��@�tX�629y�����6�xQ	�/MsSf>=�o��>J�� I�'{��)�[W>�`��,׆������I�g���q�B�����<�搅j�Ԇ�Ά�Y����e��d���n���⎼�?'6��°������1���҄"8�cb(3�������'K%p�$������y6).�z��X�ያZ����m�	l��r�6<2��Ap��[z�s'ؼ���V�`�i����CX>��[�e��:Y����Ųg���]��[���0�j�9��70лG߫E��w����J���Kq!��)[8Z��fSSӏ�E�2X3�R�ȃ*��(P"ßlfƛ5vw��W񓡠��`:Q��0>6��$v���3a�9% ݤӨµ���Kr\��;��&''H@@��ho_^¨��a���y�j�˚���]KÙ틋��nm--�/�x�I����V��.�jkk��dz�0:�8���y�z������狋�0��U�}99b�:No�zѻ����\��~
�	�ˇ;7�n�=�@�Q�r����s�䏾|7�����ۘC����߫&!I������p���+�����m�}}W���΅����~��"+���	�ުW��� =���σ*.��yꕰ��Q�zm/y���T<����������k�8\�����������v]�;Zdp���A������!���Ck��|�@YO	��jk�G�n���E��Ml2����ꉈ����tu��[qBJpgu�>Z||F�� ��m���8νB�����ghhh��U������h��w2a^�1�==�&>����ӾXﶿ2S�!n发x���Y��ϒ�o������m�!����ϕ1�t�\����e��Ʌ���湙��������db"�..������H\c������f�y�����7�ce�k������"��'̪%mil�~��5`����O���($��ym�@�|��(�wu�	W�+)Qd@?=ܜ���vs������Z^��)3��`��1h�R
׀��I�a��G_m�[H����َ�'�2ZZj�΢�}�����5#2[��[r��(�ߞ���z��,�Ej
42������xd$oJL���j|G5��Rd�O��^)4%3Sx|潥eQw���T��bWƐP20�+(��E����[��U��b�����v�.���d7����ɿa��k	�ޙ|��bU��f�%`�vEM͂<;I����m(;�����_��+i����cc�V�HCn�!yu������<0 [���@ꯖ�}���g�8N�|655����0u_�g��E�|s�5����}ު��	u��G��>�*k�	t��j�C��a�ī��l�v��s ���a!��<;�
,8ˆu�W��uD�:T������V�l�4�nna���>*zts+������C�^�ź�Wv�`�xDē/��c5i��˓�����h4av�S��D�b��Hk�Ռ�t8Yj���St������A����-'��M�,1w����f!�Ғ�������������rr�K�����<x��LS��Lx&66vHH��| ���em���	h��Y���������@c��N����B�b� /� �3۴d����o�7g���89)k�*���#���Q*���W��ц����e|�W�Ҝ�����[Z~���8�a�Tٮ[ ����$�{[��w"��ͭ��c_T��;�̸8|`����O�q?~V����۷oaFW��(��{�={�-м��gfjO��r:���?5�_Ŗ��H�T�Y�_c_�W�.��F]�4�;5��wT�B%��n]�響7�ϊ��� 0��8�*>acc�4b�ʑ�]�+,|���4N>�����~��c��3w�[�x4	��ؘr����~���p�Ƃ�Œ�O�mM�D���O�����_�.�ј
[TO휞�8��$&zw-2O�y�߽��_���#��=7�Tr���h�����m�n��ƾNRD�ĭ�Ն������RQQ�.t?7�Y��l/5��{`w�[���x,Ӓ�+��L��� ��*�;��ݸ=��ܲn�Ug���jq:�L'ATl�?cr��u�8��H��Kz{R\\�N�R~_{���ȡ�>`Y*���R���N�p�O]?!���Y=��������މ9�1Y������������ª��@���Y�Ѫ�t�,���K�D\�օ�9�x&^� `u������{+11q�ۡ���B_���ҿ�<���Ki b�z՚6vv��~����.p�������u�C�\��[��?�d��Lؐ(z�o�_�D��߹�֚��|������w�{����Pe����c�7K����a�'��P�6�
����S��"�H����Ɂa�+~��fc~��7i��8��|�v�G��/�����30��_�i��k�>$2���'��g�Y����oED����*�g�J�{O�[{8fh�Ӂ��Q{�fdd��-�*��񪥥e����<>.��	��-�AO������C._.����BK���$���@ ^�
�?���CFq�ǜʏ�B%���yyX�Z�4� P��M�乁%(���m�U��V\\�gp���=�QOw��b���۷7�]v^���Q�����c��g�j}8=����G�H�ZhXXjU����>	\��4w@�c�UX{����5ū�H�>���>���عw��߅�p��EKK���,C�;( |Ӈ��5���zmgӥ^t�WhQ��=����s�1��ˠ/�̇��ǳH��7���)鍾��f�A@������>���He���Jv��vDD�(O�9@(4�6N�m�*�[�^G�|���jhh��V�f�G�$���Zl�"�.\rA���YZu�\�ӄ=-%9�. ݏ�+,�'����q����FƠ��~~�Ix�g�V�<�Ę>aZ���q��W"v{2KKK���uEe�ySR���)q���s]��	:]"���$?~�?\����)'�gM�Rc8u�CB��׫ z�J�l��B@��� I�OHhN��Q�oaq�%���9����,��1F��������;,l-�1�[h2��Y�X����6~(1n�o��d$� �
�-�LLL����X�Mă��B6T�3�� Y�'�+���)���G��f���v/ׯ�ZINV�{^Yӵ���)������4�E��w�ZW��F^Q�b�zv:�3�tIT�<���I��oeeCN��u��|g��4�C[c�f���_�vw��To}�(�Te�7?;*�� F��Ya�nRLۿ\[r�"���E+pبE�c�y]T_��~��S�j�߽�	)i1�oC���߾��
��核���~K1W��&p%��T�ta����Y�8Ϧ�����2�C(ܞ,����=��ꐄ�Ӣ�{�~&�t��S���ԇ�ۊ3vt��a��?~�}��n���� ���铨����h"d��LIE��1@E�Yx:;��G_K�����&�}+VXc�G�C��$�l"�ȹ֪�*��+4����f�ے��#�()C.͋�w*�\�#��c��d�(����|���(��C��z��Ӯz�!G��k��,i�z��U�]*]]���Y��i��)���U�5���;��j��땽X��p�H7��ם�vv��M���J'6!�V|R�yёb��N_�|$O%-�]���r����qĐ'a{{{�"??1���.�r��l
���S�aӇ�w%2g��ȏ�Z����s���D��&9�[p���f����_�<��X��.m�,��؊C���)���Hz(�bUt<44D�K׉>@/0��7%���ؘ�g@Y���oť��
����R5Ά��LV���4�`�B�E���#��idѯ�����t����̰Y������Eke�Z�:*�_�z�B@@˖@�� _����V�'��t@!��>`V�I= 2�����O�aj�R<ؕ��Y�ݡj���i��6�`!�z~�s1.>>rX��*c�H�����D��zC�����ph��TNZ�tp�-vF�%:���:��C��N����[HGӱ�w*�)�v�P��-���񊃺���C*
�	�RR:���8y�т�id�?�.��MC���*�-�!���l�VI���cc�y�H����� �88б��͙x��bG?�nw�mmm���Vz�t\��P�(��k����ʿ��[E�%��[�F�EEVTp�Eb�Y=����$��7��R�R��%��63����R�SU��&np5��*�?&�յɒNVTT�5L��eg� ����������7Hn��u��SkP����Qվ_3����^}��V���5����րhӮ:�V���J�GDFRab�ZRRB��Ϧ ����l��RϛUU�z�-�'�,{�����>BJ^^^��/�����+���x30z8�]_�^׬o�ϣ�7�H;f��
�ц�\���H;ijXa������/}�q�7���i������`�C��B��g%õ�kj�/���)3e'�n��s{���Qd��[I	�oJ�Є����s���@�l"<<�������`��R?_]߲Uᦞ�[	<�YYY"�܊�����W�[�Q�^_�����/V���c{�ӳ� Jm�a&�}�&P�ɐ�h��.d�0�i�y��oa0l���"�L�<5���̅"���߿�ͭ�Թ��}�����*�tާI������͕�>,9
"ac��;G3a'0��d�n����Iv�)E�`�n���5R@���{�S��N��Sgܿ>�ջZ��
傸�O-4vwK�~����	|Z�d���H�ܺ��b&+m�`5����z]!��^8R?�����S�١kq�D��r�~~����nU����������	�~�W���նOO�c*��c&O�(�۹A��c�Ob<N�_QP�}�Le�%���j�I���p�E�opPp��yy�Đ�-3� %���ZDM-���uu�)������`��8!!�v�](ث�����Ս�������A��<Z��WddP�ʹ�):�J�Ɔ�����iD���I�Q�ۓ^/�n���&He���������Bϴ��/_�?6�g�ޛw����ut"�)L����.K���3�t����0P�m;;��l����������	߬��8x�[�}�{�i`S-8	�����&,,LוK�_��!���%pAb�"��Ќ\��P3��Q�>������m�W�f�RT��wt�(I�zrs�5ȅ`�� �����y�[�臙kXT�ך^h�B������f��O�5��f��_�|��U�_���IoS۲�TmVny�"{�D�	�|�H�	h�"��'s�w|E�cq&%_NڼJ�C� X6�����H92��i��|��4u�L�
H���Sf��,8�f�Y�H��5+��UV����<�'p@ �~�y�ː�͚]w�Lje$%%�2�5�k�����j휝y��-rF�����Ko"OhTy)	�ۥ�|��h�ȾZ����z�����nS5=#㣃g��S�k��f{�s��H�ՓB�;�Q�-���b�� �Cݠ��o,� ����ǻ��T�B�����}���}�
z��h��S���̝N��Y�3�$����?Q�X��\q�����3�JPRSc߫�
R�UD_[Y�؍��:1o�|�,f�
�	oJ�&u����\X���D���X���M��EѪ���Nf8���d`X�A����עEE&$~4��[��Ԥ�w0Z��0��Yo<͆�:�ơ����������i~���IH��h�]'���#�K������HBE)DI���}I![�!*$�Ⱦ�J�J��HdK3�eKB��A��,c���X������9��1�<Ͻ���~��Ͻ[����H*(� ;0�:y\�f魊yG�>(��1^K�}�8Ud��������&���G*�"�־_�kQ��ťg{�]o[�Z���j�R&3��'xP!���GaC�������\ k�dM��T����K@Ύ9�=v��
�"�"P"A
�D%9���T݀ceuZjX�� I� �s͖+��x$�} ]���O�*���R�,�^|��>����\x����F��v�dD>l@�x��{D����TK��]��W��gμbu�t )��u��a���.�!<�������Q �����e���U�4�hgg�嶽m�jҧҽt�\�ϸc�ؠL�B_>�cŦe��<�����\J��"����lWA���D�g�9	�K��׿�L����#�AG��Xr'�~�p�k�.|��!`IyucJN��^�4??m7�&B#p�l i47\�%ƴ�)�0f��m�'g%�x��	���TM3s��j�d���a���y�����c�m�~�2�i��H)�t�}17��/��@�ҝ�l���p�%(<���GK�.-}�v�O������Q�6���K��94�[��}�@Z�&��Uz����~jT�/AY������7L$��k��1(���A��¹Ӥ� ۱�x���Ya&zzz?���i���Y-�Ƨ����X���I0ۿ�n��,���w�gCmCC���ڼO���^!B�
÷S"�	�sXVruQ�`��[Z��z@E Ai?j����?��C-b�B#-!��cM�$�L<��<���YNi�o��������RWW�/%��'~`\U����ᤳ9~KYm�"��G�Pl���	�۟���%Y��[�/�v8�|�:�U0l���}���-I�z{!�h(�� ��K��G~=x��e�����|�(C�Br��F�>��f�Y,h��ݻw������\{��'��	 �ψeG�%_U���&���=ʖ�v��hS��91�{1[���)N�kу*+@��1j �T�O����~k�0=�,l�Ɲ1���8��\v1�>���#�����V�f����V�*? 4��|.�0�����������_���@$abj*�����s+y����Vg��bpu�,C�5%���7 *|}�u�ѕw6IIIO�O��>n�M�0j����W@R��~OOGh+�<y�E��x�U|���[-��*�(م&����I�{4���y����ϭ�Cy��t*�3q��4���C�&M�����c^gps/55pл�@�t`l�Xew��X��~�o2�j���Q{����w�T�:;u����.���i�X0\�TH8N�z��P����|��ȈEG�ṭ�QS�b]�'���=%a��v �M���t=K/��/�}�Ya~_1���f�Ӱ�B���*u�^����(2�e�og�'$�_���,-��F��D�\STl,|�OWWw	n�����77|!�'�3 �)����z�YYg�s81���u�%=����ro���������.Hy��&j�̜�_o%4�щYY�ihh��HI�_�yTMQ��R�f����؟L {�Y�e�����qG3|o�ͥ���s��o�{����0�����<y��#�&Z�ZF\+��W����0�{��F���'u�p
D�Y5	`Tw���6������mUD����6��G$���rۀ������������x2ݢP���3 0�|q�f�m�H-�f�>瓀ѼZ<n�*I��ޛ'L��O��/pF�{[�j�hT۔�J���چ�ec�\N��]�=9ٚ��v������ϊO7��=�����s�N����(\SWʅ�X���a a�[c��E+����֏���K1*kk�=�얺��,�Hc��a5;��1���p��]:3���'����Ǉt�������0m��7~X�-�&hq�r��J�k� ��=Sڟ�W�b<]WJ���kZq:� i��Yb��������	���ts�ΝT����^��Z����x~9e��/��ݏ�n�{ɯP3��j�uqZ��Zö��G_��+�?��6�؊���J�8q�y�\����ң�6g����[}vI�s�Qǜ�A��#yyyQ�7���srr>��sqq�������kY'h9�A�paxd��G5��0���>����Ʋ��\��$�	@�OL�����>�;\>�08����6̄5�J
x
��/>d�/[��Mj����v�AF�!�;�рlt�Q+���h���2w<�t�{|椡��Ԃ�ti��F���ꙻw�ۼ����Ox~�v�ti�������,�����ه���/��x4��ԩS�GG#q%�ʜ<�7 c;+&��r쟐�$�r*�C���0B�e9�k�,@UTL	K�E�R�9�<�X�,^���M���!,e�+ڙ,,|���!�=|��>�f�`tf��d{U���2��0�@�3µ�U��U�em�j���<0g�V�E������Bn�Kh��<y80p�k͓l*�	~��eV����=_<������E��6K���9�&E�m�=E9�cwۓ}sE��%/����cA��_�q~E!��ݞ��	����<w�L��r_:[�G��3#��d7�Z7���������x�ۚ+� ��wR�~����V��V�^{z�_6l��h��!kJ���{������5k�]�_%}��x�G������P�o{oo�����������������^�]�~�����X!{.�<|4:w�Y���;��6��eddh���ʬ[OA�$'�u����4�aZ���\{l�1���&-����jkυ+�v�)�=.z�j�`�>��.�<�&g�5���V�ʐc�/[�^ �����>.x�� c������KsT?ω��?~��85 <P o ���UN�:�a^\W�>w/n��0N��)���{��o����B�,V��E[+��}J�':s5Ɵ��}�h��D���g���n�����������be�O94D���''��zF+sVTU��p�Hk=��4t���wq[s8�"��"���vɒ�P(������s,�NW|�����I҂�*wQM�p|�+��ҋn���U�d��f�N�z6�� fǅϝ; ��]�v��eҦ�&!���@����.�?c2則�:�Uق5�� �0�kE�xu�_TUR*�ʳ�uS�����(^�����y!��C\B"?���ʪ2֩������7��ʣ����!��D�2xV]��,���a�ޏ�3�_���q �v���|+Txʼݞ�*#)�1�[�=�@���.!P �=�y����܏nN�+)Јڼ׮]��*��w�i-C��G: 2',,���.��
0���³��w뢄��g$QQQ�>�JH�oH��E}���Y�_h?�ϯ��#kn�z�����f9m�Oe���g��^��|��]���	)@���2fZ���!,,|����.�!�С�Pji�+l�_��!N.�&7�@��}!~z�.纑}�9�{)8p�Zɖ���%E�to�8�31�����X�Z��������w�qe�οb���6&�Y527���xJ9䬻մ&��3CX���K���t54ZrA6��������E��9U�T�]��'�v[�-��ٳ$���mL�\��>�Ӆ�����;9	���X�JHJ�v�3���������(ra�_M!c�
W��q�~~R^�������ڂ����,C�[Y�Rl�|y��������S*�w�-j��ocnEOB}��zI񌚚���i>>Ǯw�DD:���ޞ��@��钵���c���������S�u��z���w���@Є�t�'��캟
0���U�j5xL����*,V}�W\��hK/���ޫ+ng���&� T���:�1ϓjzzLų�6
%q}��~�K�
�t�_`�e�Jq�UutÀ�h"�>m�]*��@:���}��1 �j�?B�+d~��@�|�ﯮ�13P�?��j��˗/���jkkw;�3���_�EL+r�3���{����e�3��Ƕ���ulK�@

��
��>��ǘ�gvz}j�ţt�șQ5/�o�QH�v;
Jʁ�er{��gT��\'O��]@�KX�q���͹�tfW��s�o�w(G6�Wq����E�&F��	�	��`������9���]�.� v Vx􀂋
u,x��y�u�_?{M+W��Y�E*6�����<�_���t��w6����o�~~:MM�.�ɟ���Jw;�gc%sš5���0E���7&�M%�.���0_�Q��~��^��)%�S�<�&7���0�L}�4�h,���p	s�?唴F�����L���^������؞�/;���?j5�W����l���Y�y��E�;?��;U����cOrs��`���ԔT'!WuU��Ky�*��V��
d��g�D�Ǥ�0��W�@}�PU-�n{*m�P���*^�����v�@*?������P&��W�i/[2��+���^�p8�?քq	��gV�g�ՙ��dy�?i3�]���Kְ�7�`�XҜ�0:>f���@
Юj�A&te�չ�(�og��T����+�q�*_��(!{%�1��>�_1�Y�[����m�y���0ǲ ���~J���/x�͋�o��n��Xvx��S�H�恵�3d�DFF��|�[mm6���й����z�A��5��o%ߏMH`��+b��Nb��>/:P�#	�����R}���G]b23;� H1]��H�w��jϣI(�~7��g%>�����"���[
7�QPU�ZZ¼X�m�l���ʘt,hll���ѯ3�~�3��yi���8�v�|R[|h�i��h�XI'8�� ����pb���%w*��xm�EcfVVr::�UUU���g���;:ntX��Up����Q�x0�3yj$�-3�����I����ܣ�>W^�;F���^.՘�^^21�\�߿�WStc�k�LM9�3������f���.7�u��YVL�:�q�� h{�B�!	R"�<9�焅�"����i\ɺ����z�g�"o���w|z����Yҵyዕ|�_�d ŋ�W�,��@v����=�ϗ�#��F�TO�<��ϼ+�C\'�hr�Y	��@ �簬LO��H���{ܴ�ѵqfu55:�#rw�j,��:��u�[y��e��wz�:�rFW��R$1=}_f�z�|�l��_@[?^UQ	&,����S�u�t�C�߿� 4��˶+�����{]O/ XX)���<�4�����l�H��@��X)�/���6���4^�:���Ǐ?\�b�V�ʮ[�H�g��i?mu^�Tj=�����#���#�U�E�LsO��2����ms�;{>�ԥ(�LF�#y�4|�f��Ӵ�jb�����p�8�f��g ��k����U7)�a/��WVQ�I��"##�|�sH�C@m����_�2�hii�6ǯ̡�ZYY���OA<�=�<�ʎ����*MM��QQ��|�ǥ7�sssG2#������{����G��989�yx����.ik��ͅ�*���ω򡧩1̗��M��a��-���䳬Sh���hya詫�gw���q)2(���a��,�����~�r���Gβ���*?�oZ��pD
�*���8����G@Vu�UUW��ퟛ����]���D�	�:�Z[[��������_��� vm�G�,r\X��ɓ'����E�P��oT�Q&���e�Ԥ28�	�+bӗ��*����	��w`�L���aA󨬓�CrJ�|�����i `@aR>wK����V�ge�--fL�кM}��V�nkӮ� VucM��'O�)����{�=���PW�2�ʫE�������<l�w�o�J�;��ĳ�P�*�3}m֟;J
�c�����g^�A���|�۷���P�?��F����;
����@�壘iX�c,���e��w�L�l�{��&|ˋvk5��;����@>NO<]ǹ��I ��	`<i3�Kp��tG@�4453W΁�u����B���C���lY��3XYY}����NSaP���Y�QJs�_XPL�����J�렽��ϯZ�~7{�>�L�#���9��Ƙ?<;T��_���m��+"PS�o39R�žٜ�{����s��o.��H~	ǒ7*�����|�?��F������[0V�B˭��Û�D1���(G�6H��:/��#sp��vC��B����O�5���T�.�64d<�q�����\��.��+�'�R�͢�,{�}P�@�^R"?�#�'�	��r��<HZ8j�����5�%$D/_*L߹OGCC�mL> (�����S�#��^�d�C>3Ķq�ʕ+M��h:ii�q�ǵ���r$@k�*?�	$��W��=�s��2:���]G�H� \�l�b�~a��8X'گ�K!���QO���l^��B��F����e�֠DUo�d�ט��ʺ�����[M�������,��&��n�`�ٳ�K̭��*�5�GK˻tO�$@��O9����_�<��EX��^P��2�x��9uި?@>/��@��2c��ش[��F��i��P�j�Э���d��~&7����2?/�aj�z�xs-1g2��
o7��o�.|��9�w�ͯ�.hܺ�QKխ=����7��4a_v�K_	
pwϡJFC��+nn��us�cb*>�*0�|���n�3�O��v*������4@�Ù��������#��s.��9.�gÎ;��~���'.�:|w��b+b�+���އ��Z�2�?0�u��>&#���l(w���V�|��Դ���߃rVt�`����?f4��KA�|�jc"���%�3�\\���+@��`���+̧J�2�l��\�g4���)UR�?�4̗�R�KCf��/5��tt������?��n=C���"�D/ʪ?�$�p5@_$� ��v���۷o/�k˧;�_XA���������/�ٝ���|�*�*��u�
�,��;n��O�&�n���A������f��mH.j)���M��802tO�|7鮵�d�ர�@.���T_�B����@f����U���)�,W�"��D&�_p����)aָ	_�봼�94��]p�ma�U�p��L���D�������l�E:���� B�����~AA���g�����1�/�@���=Y;3�åY˥~�jd e&9ޓ	T!T����١% \�R��^�)g[�rHc5�[���P�a�=�0A9�#_c���ԇ+�o�nK�o���^�B	9YAB%�a����"~�'��ɮL9�6�#����^�{�Z2���N��w�du<K� @��;��f�6�k�����`��`%\��@��%&&.�������2���i�I�g���3<<�����H�� pk�1�w�.8�A��v�����f;��)ff|���AL�w�×/�V~'J��ޗY�g��j����a� ~xN�� �]�hiQ־�j�N�'��0�!�']n#�o�~�9�h��I� gO�P�,��up������;9�e_��}�̤��oO�8�j$������2�9MM���6�ŉ/�@�.�;�����XX\|������Tn��j�	�3��>� ������A"Z�Ū�H����V��U����c��Y�X�f������ՖTx��CPa��kG���+H�V���f}��̙3��Ƿ`O�e�]!��|�k�n@@�~f�tO�^\\�ZC�Q\��^�"��-��<"9C�ߓ������=H���{t���4p��>ѲfP&A�-YV���� ���Y�^���p��EX�!�w}��6�#�~p�cT��)8ݗ4�(.,,�<SF	ߩFI�ͥ7\��ʚ<�\��}����1Q�N� Q_:�*��K��Kx֨Jiae�ت�@���C1�ݫ���O���jj]�&.Q���[5�-���0�d�N�j�D��į�sMtd_Q���<)c�d�8TAYYK�$'�@���]���}}!�V%�hfW5� JW���!8@�g���z��lt��0�>	!�6��0RN-P��΃�����Gf��U!{{��_�EEEK8�'��D��It?����k J�'����� ��cu��:�ck-��h�/ )��~���j5��a䊃�0ܗ���!X膇�4a)dژ��/;d�T@��Yv�YvϺ�w;#qdss����1 k���g�����R�`���e�~i�kJ�`JhN�T����P�4�Q��ccc3et���(�i�'�2 �Aǡ������4�@�������1���{ϟ?���r�8�#Ϣ�a��օ�19%%��������j��@k�y,��!��P�#qn�@(J\X���м ��w��B�, �;w�\v���u	�/\�0d<������1Pw褊�%�>�U�5�:��AV�%o0���p߷��MY�|�h��=�B��&�"�:�:.��훋��>������|�8�0�)H�W--�w�BQ�6^٭����>�hn��+.u�[kk�7�)]]����/(x�¥Q94�$­[��Ӡ"��i^�<�מe;t�eDD"�I@������[� �=�ܾ��?���\<�MFI�-�!��0��=�{�
�����ߺ�� P�O>�����oT��k��3�h�쁝������*n����wc�����H�q,qnS��7Ѵ�kw|�O����}�]�|��0�)��#�y\�W1s�H��H1HR9��>O���W�z�ܞ#�i&a<�[tDF�L�"`��/�I���F88���.}��ȑW�12�Q��D���GP�&ϭm8H�9z��Ǐ�p�CJ*(�^�{���7� �"$*����Q5���L�ЇI-;�v-//q��_H�ȠQQQ�;#���}�8���|�:Zji��+��Pʲ7���O��TUi��i1`_X�����
 .&��x
Oɖ~\>�����Χ�`��KJJ��SM����0���(���~���ӟ��1R.I���][s�{�W�t��;��X_�������̽�@��# ����E��o���Ha�EY��Հ�ze55j]��]N��i�El�jR������&*4V�&z���Gt�6F��t�Q��ACG8��<�;~������Od��9.�f]��.�����=Tr
{��z��`�9xy���Ϟ�&�qd	�]b�<gѠ��+� ^R��?*�p��P�� `ܠ%==n]`z�k<�u}jz�|̷��W� 8Pcc㗆Lр�!��>��x���^F[S�������%s���W������I��i�T�N-@�s��k��k�'���x~ʩڭo.�W�Lf�W������A\��M�˕/ k�<��mR��(�_�X�hX��}��.Z����Y1�9��p�A���;��q�����?�J6����3ebv�ʅs����ˮBL�������<Z1ȁ�12^�W��yU/5E3�#��+��gMeu���82�C��ԩp��l�S�����	@�:����+��gi��1p9U/S�^�u��o6�ƃV���l���[Ӯ:1�n��}�*S5�[R5m��������-��
���������|�+�ԡ<|�����[��.'F��B�[^Fbn��r�Z4�]Lc�4~��Z���Ļ�h��zD�E����gd�^܈����7���V灷@��Wgf�<#97��2���Y$�P�������ϊ��@�Õ��@6��������mv�}�D�kQ_��:H:�Z��g�v�WQow��N��C���_x޹P��K�g��I"Vr�6�ռh����	��o�����LpwsI}}}l��x�T��6����`�٥���|���ttC@�ڎ�et�0��I�L�0�0p=��<j?X�:���*��X�1B�6鸪��y�����#���s�E��P@���"��j������}��0R��w���,n�����AQ~��8ш�w�]�8��p�s� 򈛛[�,M�����ڇ��Ѝx<���1?�/�Pv�jj|K��H��	>pi���	j�hc�x����W��t=6�R]�6O&3ŕˬ�SK�6].=}��f�gՂ-S?��x���c mO�����8МR�h��nD�3����{�N#�{{U��|�����Y�`[~Φۡ_�I��䟐��S������r��Z�&� 3�pA�{3t7u/�s����X�nƹ�	�qKnVL��$�ɗ����>� �-_�IA#��i�^��T�뙓RL��#�E�2�zf^����`ߗ&���(�)�ͣc����p��U�팎p��q���n�&��ϼ�w-�~!NJ<��{4O/�yc��$k.�u,u���|Fg�pD6[�þ+�i��HP$��gD/���Iە��Ǳ\еX�q�WJgf��=:��n�&�S�,�w��Nac����|�@ ��G��~������K����w������c Cvo� $~�s��] ��> y������8�4��%��lF�{\)]E9�L!���B�.�*.���t���4G��d��Q��x�z�+����{�v�R�S��`��}�2ە����G`�ϗ�ӵ�q0�b��/�i�·�UKQ����%��q��h?
Ȱ��XI'�o9�.����ÙX���Oqy!.�α(?��)П~�A�!�iN��3bU�jX�7{>5	��pm^mc�K}�4��D6�i$$s����6[�GG��۬_�'�d��hB暅���L]����g:c�>Qc@�#�*��*.7�Mo�O�C����j1�i+� �����q���Ƃ!�=���	d|�~�fZn������'�D;!�\⪫e�g;PK� ��o^|�d���T7�X��w�qd|�����Vs����ww}�Gn���Gw�}�:[�+���5h��	m���	%��g5H�|�� `����7O�c��:�5�����K���ܬ�㩡��2���-yE���/}Vn���ي�&7�Ll%�%�tR3��p��0ަQO��vX��B3��yr�O��-��
���U��ǁ�P�d���W��*4��݉�����h�a* �+־7T�ɬ,�R^؟�=�����/1���i~�ZslH,��G1a@mᰳ�lC�O��8z��k�q�ϯZ�_�^a �cae���|�ž��@=�g������7�0X<DHS+�`����E��	���ч{�J������!����9���徻��|��<ѰBڠ��;^�lہ�%����Xh#<�v��I%�!��}�y/z��j��VSY��_�oPx�pm�q��Ѐ=]�����\��
��5p��;�9$���q0e��ȧ���]X
���[M~g�?�d+�����A��(nu��-�>W1��̺�#���0ϒ�=����Mg;�B=p�k�6��TML��y�$F"p���E��O4���Į���'�Ty�������Y��P��_�祎����o�1�{����F��}�G�*�֜����`/$rR|�<��|:���?�Jxm�^�7��ro�.���m*�����ڿ�~`�U������T�$^Sx)�'x=���� ��_�p��:ޞ)�z�m��S�UϽ��7C��֯=�������.З�X��.��c٩C�C��@���c{r}%sC�_��A�L'��_l���6^�n�>e?w?v��O��
I9�.���ݭ"X]�E(�$
��㕌�3��zF.0RRR�C+g�P&��n�AߟC6@�j2��"�<�y/>��^+<[��2'F��ŊY/��~�O�o+s�����m�w�w"���g8��&�ap@�L��W���v#��M&3F$%%���Fr䷮�h\��eo����PH��G����$$9$���j�5a\�Q��'��Yt>����*	/х�F��"$��g�����$(�9���6��	�dA ���{q���� ���;ĥd�f��ӧO샋\�83��d�Ɉ��&�,-�X��ʌ��OMM]�p���-�=�I���zՐ���t���zN&a���F=��Ң^k�HM���kB�4�,�d����
�h~
��Tm8C��~ƕ7F�SM3V��%��Jį}K�u����x�F��c$��8�+w�"R���P_����󵶓oq�Bx��n◐ݩ���0���������h;�g����4R ����Z�4e�����-GY0Y��g�0QV��ݿU�ЧowV�nm�U
�t����0�@�Hw�h��4*���\Q�ǵ0���=^����B<��`�ܹ!,{�*{{4����w�g��6���iN)1p8w�߽(j�*�C��G��tp�=�o��G%��g)��x荺�4��(�U�C��7ݪ�?���8�PW�	�~?�쐉�j[����DK��#�`�ma��F�� Jy:;c&x/&Z��)��P����O[]�Mt��n3�[�AW��a�
z9���~�;��
����nn��9����OP��Y7C� ���=�p{����ؒ==#Z�&/�k{	�s�k���&�*��n�/��)�O���TI���L����D*��0��%��3�L,>�iAZ2�Y�h� ��`N��\�Lv���=ݓ�/���'0����:E����K���<3���·���_�y*����'��b���o����x�����"��Nz5����#�5�IqR���{OvO5�˨y�]�Z4A�Ҟ3�QWh1�n�$�m�����+��ب�r��Li����
�ui��x�hg�+%��q<	�Z�Q²��
��PT����.��!L��g��&[q7T�p�r�S��Y�pq �y枒�����G��$�f�0��Ս�>V=aQz���W4S�[��`Z�A��&�Z�-=M������ &A�LM:J�ĸ�t�3V����2�y9�jr2ջ��E��.L�<K���3:�1��ggo޼y�)8��Y�С�� �!��=�{A(�<��J� tE��Fg!ŵ~PR�}��?��s.������xi(�5�n�0E �X��17w�zNv�9<f������.Vg� V�舷�Rg8_r�z�gl��u�K�}=\a�p<hN�^[��UR�"������z4-mB�Lk�n{�}���o�R�կxu���l�����(u@]���y�MV��+�g\�p(a��Ǯ��7���؏�eMH��x�4�z�`�W�5��Wv�.)�i�g�x�q���
~�SƖ�p�NߖR5ۇ6��yϱ��z^���*��_�?QgjM���|�x�f�E�%Ц(�8}Vc � ���#@TZ��{���ZM��aK��u}b�T8��yer��Ӟ��<^\V�o���6�us�`(q���ď�Z*�~���/
��W�e�5�8�����ae�����ط82���9���V�C�c��]a��hj��'�N�(�GE���-�ˠc�o��U��L%y?9�iƎ}�����OA!1��$��Ky��YEP�dY�O	�������%��/��'%�^9�{bf��I���3'��p��Ӂ�p�\iO7��2�?���UXfKe��{�Q��o�0YWq⭙{�~�yrax2�ӟ�ЫҢ'���N/���|�Q������	�~ �R�M��)���T=
�*Ĵ��l�ܕ��%>�+X�ŉNI�8R�u7F@�����gDkRɧ5�����Ԛ���$�8�M�;M#*����\���3Ut_��/�L�w-�;6�8�T���}$	�fek��Ь���8�?�c-��x�C vq��̷|�v��a�'&*@�������	 �(G>vO�A���}����� ��5y�Z`�6�1kZ�Ie���d6��JS�rs��)d��[��
n����>nSS}I�ˎaD}�hRE0H/|�Gˉ�"l�}�haj���r:KV�q&L2��[�~�;bn�H�͆����S����cگ�bN����1����ƾ�,�9V���_N�:�fq��5rH���ٔ�Ő}��5(ϧ�w�	:��U�>><{z,:�K���O��2�Z��H���͊a���_PB�V�O 3/mkBh��ڦ	d�������d����/�h*��A����}׵'�>������*io���"�Gh�α�Z4�GwSY�/���?t�.��؉kٕ��q�eTz�JĪ���V�o)�EC��a����=�*�; ���:bY�a���J--�0!;��#C|�@)�gi)�wd w�z���[W�G�Zu��R���Er�O��ʻ[�Lp��a@*�1�tB�ǝg
��_��u�TӣQݤ:�)p��|b�e��/r�؄���8��B���ﻘ����41]���QQʜ�\���tA�7�ʗ�
B�<b ��a$�~��;Ͱ}s������ ހ4��8��<lq
q������\��7�`!�HS�1������O��l�2����e��`@��r�
�PL:�/n���C�.��!�a)�wE�c>FeO�Iٝ�����V���jv�h�P�BJwpYD�Ѫ��23)�H���#6��V�rÝ,��}�).��ʗ0�pOSC��k��W�{n|�m��,p/A9��$��y��Y�2�\ߋ���ݶ)r�%�������0��tB�E�Uhzܠ���c���J��x���)0{��3��(T@��G����h�p2#�Jz�R�9�{�:w�ʙ�Z�u�%'f'`��p�N@��Պۉ��Fg��8u���;�g^��SP��� �}��9����\�X��nHu{�BP�A��_-�.������f9|�%�3��v��f�ʆo��N�nXy���
nop�`dR,��vdC_�8`�5��muFg�Z��u��ǖ���#�Ǫ��>�$�� �^VV��y6bҊ�\Zr���%��{�VV�V+���?�-���Ufզ�
��܇�ɐ�~�-����hf��z�C�l�Ä1�zNJ (|�{�z2�"�]�TvNĤ���*��Q�)�w����H���8cA�$�o�]vǍ�m�����{����������m��u�˦!�J���m�ihHe���]:�,W��I�X�Ҫ�:Ź@���.��Ri�武�3��(��7O���|m7&Fy\i>��&Y3�D����v��4(�������~��˒�Ǎ�W�s|�n�{�^e;�9ѵ5�TO���J�;��S�Y��lt��_�yq�𾛛��:S�U�H�Gn����KG�=R�+��`M��fjH��RįTz���pN�v�{s�L�2۶�L
�b��#{�v����K�q(�������/�zڷǧ�\}\��K��c��\��\f�(;Tu��I�Te�Ɛ5�pe�3��{�p8��u�v�^��A��&��� �C}ĢI�e�q{���y���ussNeL�<�otks��?ei�]���=X�f9����g��(��� 0�!��8,�z��K`'�؃�g��dR��6�^<	��F-,�^ P�����4U7�؟�(����n9��)����,��^a5��?%�AM�4(v�@Uk�9�.��-�*+j5?inT}���$�܁�F3�<�kh-�5�=�3��z�I��vʭ�4�j�?�,ǎ�mߙ�b;�E�_�j)>�NF��%[������V��3m_ěj2��cS?�B�Ǥ��B�n*���хU���j�D�SX�)`8k�ɨ(���%����<H	� Ս� �vl��!Tt��{C���Q��0�����@ɾV�l4ou+��ڃ�'��,�ՀC�i���� �e
N�������B�Ċ=�Wb⬆V����Q����q�(�ͥ��C���a�	��voOC���hp��wI��3��}N��;3���Z�"�b�3�c�.�3}s�h�ۅ�sc,#!eF�ݮ��4Z��{���u���{�mw0���`�/�Ev�S����G�E�s��L(�b���D�!L�WZ�����Z��qQw��VY	�@3u��q�����UX��g'?��5*���vOp���{R*}�G�YLB"��B�i��|U�s�e)�1(�U�T/J�� �7�Vq|����a�`���ص<_�3��&�bĠQ�/�H긐jƭ��A ��9��,�q��ߔѮ�;�7Ӥ�������qcOc�ʁ��j"w��W�N.��J��Z�����|�b]��%ѷƭd��W-�W�{���x$���M�LE9V��
)t'#u7<"ȶ��B� ��%�Ğ*�9�m{��"��D����� ��'M�`�����(� �f]rG�u8���k�5qD�EZh����I���I#��h��jȖ�����{��}��C�Ԣ!��\�I�H>�߁U=V>�#zGo����uD���ʕf�,�K�k�������"��')�"��N��kh�}�is��x�a@�ґ�ŧ)7�S�?@�voO�]_���k��(|_+���Ÿ�Dl_o���b�5��`R49֜�r�i�8�c
�@�7f����P��,���$�՚�TO�C�!U�����>>�C�3�pLV���06��0���+QE'a5��[!��H[?��~l"�i
�W��+ظ��)	����xr S��}m֟�C���N%�4t�)����m7ɳ��,�2��+l���v�;���^����!�'�Q��4S��"FzIE\�s�9z��	�]�^���ѽ�x����(U���>��.����dh��{�b�ׄ3��ee�i�"Az��J?ך�]"L��9;���k�~	,����YϠ���ɉ��,2
���߿�9�s�y�/Iϒ	ʔ��	x��t�
d<Y�~b?Y�
����؜�"$��΂��j���k�]���_�_m��vz�h�� ��Uc�j�=v��A�_c���z�$����8�>�[��ؖ#��ahV�jhE��:{k2;̈́��/�j���6��&�DR+r?r1op��S� F0�y���:����ݼy��zNZ#��M���n8qB��f�Ž>~�qh-H�_PL�ں?�*۸u2�� �����XYp����.-Z���K쵮���b�3;���~qg�@�B��wESs�na��]����5E��4��#���i�IF��ʊ�KȦGw/*c�C��wB�u��1Í���&٬���Ԛ��n����4\Z��UH�fv+bΑ���uf�2��*����5�C���z�-(�6�� t�%��ú7�Ѕ���7��lK���־�W�-T=7Iq�^�<��f���T:�%��18����]��?4������v�?�y0"��?-�8�*r>Ŷ ���k�O�"�PI��wW�F`�Vn���� �9lPAAA�c��̶��[��f'3��G7F}/)�N!a.)$Hw�j2=\c
�z�:�3L�(j?he3�hQ������j�SL�8��.��Itk� c�pδ�D���׼|��]>n����3cGzM�HOF���{�z��V��I�����!��
���I��E$�Q��i��&ZuUG���p�vcceiĤ�o�qNaO�;� �@�e���o���zevC�K��c�c�����(J���D���9��΃�ӧO/��ɵX%U�	�q��<p �Ҕ�;���7-(`�A�kۮF��X3�*yu�S��J� ���B��4�̏6ϖ�y�-��*�#�zX�#g��Ңv���_��@j���eh�4Cw���Go��Zu����$fy[|VJ�O�_��e2�v}ߣ��X�˶̍�Lº�#����o�$�~i�DM����������c�p�v��s��6T���8��O�����}CڙA�r�u��a�ZE}�DA?�ί�6�:���\���Ƽ��K���i�
�a��%�	�D��bA3ulaa&�?���]�?�i�� j�o/I�
��9&�sqB�«�ӓ8��z;h!p�.ڠ8��ߘ���B���5R"���o�����&� �P^��'v�8;E��<;��*� 8z�3tzۋ�}V��^+c[��6��~����|�����'Dq�����R
��J=Z�;���ۿ���̽7��
�JԘ�C|����n�Er�5pY'4�j���xz�J�J��*1�B���j�xiNfcn�V����D����%?��v!�� ������yD���/�!��:^:w-,xG-� Y�q��v��w�|AK��W4H�J��X�V[��uAoH�������Y��y��NS�������M�k1�Qxq��{2��w��3�t�EzK-��Ǐ�~ɰ�Ȏ�^��������js�H���ovҌ���AF�Ɛ� ��D��K_�/<�fn�����W+��d@��4��m�.~�&,�D�5�!ҭ�N u��f���Z�^�K�?R���#>|���CF}qN�8`��6:
V��N��������>|���L��j[š
��p�rs݌���{�S����Z*�D�,${D�c4HF$+[���c��d��U!d��g�s�̬#��c|�sz������_�\:������~��o�/W�0��hL�;|ԛ������0��M6�K��i��m�t+*~2|��̭(c���������^f4�u��H9镕���Y�Y�Ж���R"zL�Vrְ~����t�1���$��^Z|�i�yʭ/0�|}�۷o\S��C2؃�&�ZN���%pI��u�g�4��̤���~��4zȕ<��@O�q&�|z�j�Tf/k�n ?>����y2�~�@
N]#@Ŋv)�1|z�cت� �])��駈���n����C��B�����>���@[�"k%ZF�%[�4V�q��c_����Q(���bm���C�, ��8KJ�{�/�ɦ�^ʼ�H�rYfOa�ݕ�	��,�)�"��+F���2
��\��;�Ж��{�k<�$M�����d�	l��� �SD]R4��B��B�\�a���AC��_<#��2zTFC���������ݞ��=��������eP�L���$�t�";E*���QG���*?�kt�L�:�:�C�jB>;�T�%�RO�T��U~%��yɁ��_��,�@��G�0�c%�=��o�444&|���<A���ϯ(�4�E�]�>�y|Ǔ��Ͱ�ܕ��"�a���$�%\0+ x���`_�]!�6�D��� ��t���C�i���[Q�[��+:5k:+m5�mPzg�j墜"��Б�{Qv���	 !�_+�P�����~p]2��r$';a��)�-)���P�<�uv ���$���:O1����}��z�e7j����8��� r��+�a^£�ɘz��q����qr&�}.999����GrŻJ׶�藺ϲ�YF^V����E@�"qw#`h$k(�SSs��q�;�C<�s��r���8}���ࡷ_X;׏�uK���ޙxm5]*{`�{��d�P���U�=��j�1��Ӕ��"����d2W���VJS/��U8����Yv���^�al��� m��*OA0�m�<n�ɔ[���Z��uX4Q�"D��˝zxH�_Z��V=R�Y$��c�-LCp�VM:�'y�Bp�b4M��������ً[x@-��!H���bQ(�C
,ľ7/���1��kնj�4�V��F�it�������Ҥ����{��w���N�:���?A��+թ=+J��ar�uY��.��So+Y����v�V"��ڪ>���`�� �n�1<��pfDa�'���Q	f�kz˴d���>c=��� >^ޟ�����������:
M�N���\�|mW#�x�4AB���M{�	�ÊBO�L ���L����X�ؑ�f�.9����������g��OYc�s��h���&&&rE�	�r`jn�A��N����S-v��#���~��EEj��͚1�)�S���(k;��.wǫ���"�7_+u��\�ї��;���d��4:�>���w
1$�fy���7�`^��[�>��h[V�<��h�J�'f��)�#:�='kO񿕱�wy��$
S[�4�Z��Ɔ�ư�U.��s��VI�g��ZlĎh��+��ݛ����Б��2叽UR;umDV@�Jv���k$���I���������c?��3�( ��;�+ë���w�����-|�y��!$���骒��B���HiOB���q�X��Þr[��X���cj�ܿ��%\�&���躼��	�bWq\"�_��j�7V�v  G#7g@/�ʒZ���O���W��F��O  (��J9AP����^�G�9��(<�F��U��Ob��0���jY�#��
g�G.Wcs����|栊�ꊗ��tJI\��n$I_�5N�\���q\�h��)����ř��ܭx�І.�f�U���7���޿����/�I�S(�?����2�\x��4��j��'��XZrz�x���v����[J�������8�<cu�&�e�f�j�q���F��0��� ���ޫ��+�~��t���. ���dZ�; ����������ʺ�����&�.qJ{��S�U�#'B�@���%���`�Kb�X������'��$0����!��|�XJ�T�n޿��K�E,�ۅ��.E�H6�B��2{��n�Lno��v!e(��B�q��[".��\f�@a���Ê��\Ї5A���HL>�iIٖ����ژ�P�]^�8x�)V���_��xH(w!�`�*Qҳ|�zCfZ�}d�����%iC�@O߼]<? �6ǐ}8$���"��W�߽��JT�Ѩ.������P�9~���'�t�IP�?����x�D�\N�bu���������n��&㝂�n��{����j�΂QQQ#c;#�9cN�B�FF�ջp5|�B^��\l��1���E(2�%��`ea.`l3i,���#��W{��n�DT�2f
-<�US��o'Ϯ�{o����y��Y�Ts�u��h��h�O62f��8s�,���W�nL����	(|�w��ۂ�_�ߞ"X�=g�O�"L�<6>3��yoOb�P��@�f�'e�w�$�ĸ�/�V�9w�B��	P�`�r�0NR4#vp�g��=&�z[���܏xo}J䑊)b	TPsR�kZsb.#e���c%� �`���R�3�E���n��� X�z}w9o�[^.��Kٌ�^�$����!��&�*���Ti�����Z�|aa�1$-<J����Ў��e�������kО't���"m���7��W�,�tH�a�EGc5@G >
df�.V"r+&F���Х\:�Xs����i"3#90#ٝ���;~(���+;C!��T/̭-��uU��c8�DvI�wIb��@|�PW7��q2����������el�e<e�Cd�W]�!*ɏK>126f��Xi(�P�J ]j�Mi�̉Y�q��w�[���x�Zo+�:��w[��涫q��n���Z�����x��Ne=łc�z�6�Ҽ@�XA64�'���ߟښҸ�*��1n'B�*��E �F`f|Z˾�F�toI�Jæ���H�Պ˼�y:���S�G�a82�N��:�B��D���Kn�!��'�},Y��	���N�z';|J���-D���\��燲b�Og�N��sE��W鯓�y�٘p�o�����"?_E��v��U���v��DEF n��|�*nM>��(ʱ���i����S�i���h��!wX#�8��.�O��Ϧ���L,�;�e��7��~|��S��,�@xT�*��}C������=5��`�N�r���&�E�n��&'�f&6�l��$'-��D#5�T���͐�$*�v���.L"������S1{p�"&

�d������]�l��T�g� ��D�0A�/�.�Tt����B�v
U�JH��Dφ���:���ය�w�&�|�r��X��Y�����^��f"�2.�^A�d���/�L�0f����k��b�K+��,ty䢃y�";�2�&��j�z]6=~NJ�sʳ���;�@�Qt����h ���U���Y�<OW�F�ŭ�?�wʺ����ZS5V��3䰜�Ά]�зk��tT-�AL\Dz���%\���V0�ה��h���@*���]�G��Z�v#𓍷�������DV��uɒ���K|l�A&D�����{�N�zT��jI���OaB/t V>�!؛�Q��z;X��nk���f�/栄��(�Ԭu���crgWBK�y�0�5���㝤t!w����H`x\ܺ�o�?h��u��	+�P�*�1z�]o
�6����h��_��4XA:�w��視�6�J�����f�q�.���*w��V�����ɻ�:�(����9>=<����{�����f"�E9�����n۫��?Qמ�~ҁ,��
��M����ou�s�3)K� �y *���w�H�!v[[�s^f �nnn~��`U=^��������n�x��W�Lz�y ���P�60&ǎ쟾Iڐ�3�!�x`���c�u��Q�)3���}�J�^�/P,�œz�1�b`�w��
.�cq07���C-�� �]_� X���Ш�r�J^s����f�f[2��`�2�a~o+eP��3ޔw[�NH`��̪�NZz[3(W}|�N��V�J�Iy2ֶ	�;@.@ؚA`�顆U��4
��_�%����+���L�Dx!��A,��ѱ��ߓ��.�p]�I�{��`��*��E�/���P`0f���kb����?���#炇e'yv�� ڥ��q�8��K��z[�/��ʯ�frC7e4��	��h��>�*~��i�k�\?d�L��5�پ��b�?�h�ԩS�l}Xr<�OoK孇-�gF8��x�DA`s0�Y2�,���D��#������0#Z�r'���ؒZ&?����R�h�g��T��2$$$`��ݫ���1�p����K�a���D��дS��e�]I�w,5��t��>\ut�1��r�D`x�ݍR2�j_+�����׬Ƽg)�w� jɏ�Q䗕�O���� :���bmm�nϓ������D!�EEcp��5Z����o�4�������m,���ӳ��|`aM�a��z���m�IB�*�A1Q��{�.���WVǸ�T3t�B�u�X���U�����Z�Q�<�y0�p(O���j��?��(VP�k�� ȟcw�_�8�9��rCC-)� ��ȁ۹��OX�34�W,r�i�e�j�?��j����W;Go�6AQQ��F���>�w];�`D(s���k�%5��͵��Dn�}���&���y+��O�/rR@�`��(���#Rb�f����Z��%�4��r�*��EN���n�9kOݡ���ކ��33fE�}�ݼIJ��-��~��?�;��q �����G�"gů���S�U�HI���Z[�$܅#HvNİɥ/���	�a2f�|@�0��c6��Jz����n��{�=��4��@}'�7v��Z������ `&>����d� �E.�
��ϕ�9k2�l��L���b� 4#S�Kד�z�
2tU���kF#v�"���bw���<��_=`��%����Q��V�#�탃`K�X�L�l~A�Y2F.D��>��.�'Fz�yx>���ʻ6��D��Q���(��������p���X��M����E`*u��&Q������v�ݍ����;}�y�l-~����~���<q��'���蘘�>+�*�k{�S�- �(+��z��o"[����k��]g涽���U�XJl�������>�r*�PNDkh%SEWGG��p �	@/����ת�����?�uG�|zH|��{�	�CN�_�2������״��1���#t�۪����kD�1i�l��Ϋ���N�|:��~dąMn(�b�J���*X�- r�srs�/�Iy�I2�#\���V�V�K<Lclt �CQl9wx�Cܟć�Z��)	�=�鶔�����?������$n�t������nL4���i�aw���J߁���F��W�S�T4��b]�6�u&l�ܡ@൉����,����Jx�&���3&��?.r��D~ykIGç�����lf�ˍZ��)d�}�M��NvI�lu��A�YJY'��u%U�8��1�����������0��\� �s� �1Y*��u����3��d9��w6$^��N�m�Qv�)�%V(}�ӯ_��T����k�{K���y�d�7����~=:H�[Q[=��n�~o7���>���	���/� >��$O�7�g����"���%���M���ؔ~~n1�C�no���J�9�+�c��9� 2��|��2��:]�uCjw��D�PL+���S������IG^�(	��$��m���2�,� ������?�\D~�6��R���*��S�X����"������IA�j�����p�j$��֤u�l�i�G0<T,::X�h	�!����n���q��ڐB@!�q2O�*`����ЙM�5!jF��yl��P��2Kl� �	�x q۟L:s������w#G99Ծ�H{����I�#搦I18Z�A��55uk2>X����l�\U�@�Hk[�(����η��>j����O���Ӽ��ښ&�	����;ib޻ :5<=r<U#;J� ���_�a�]5v3�^�$� ��P2zz��e��Gq�9Xl-��������bjV��T�Fo���{9��!7�ξ?�MH�(t���W�C�nԏy���Ο5zef�uȕ�)L��U<tzzzpp����É�^�&N�4O�O�)K���%qP?��ۂ
�V����W%ӏ�� ��S�]M{;?J'��o9�*�	�0����ߟ:�� ��0����`G���c���ơ� h(�w<�><mF���P��&� J�M����Vg�d���F��������umAD* �&��~t�T��v/њ�m/�v6��M7�n�O�E�(��Qr��-).�=�T0v�N9��O�$=n�l����B^��FО��se�MAQ�ͫ��?m�a&dU�݂FC��8��6Z�h&��t_DU�g����J~qp�4^s��i����&�P������r�^�e���C�k
���c$N*i��e�~��sV�U�w�\�N��*(vv��m��?��o���	U2����������X��=3�LV[g�����M�O1՞��ս����;1�1	��8(þ]��:��4qs��ڀ���{҃[Q�GR����f|�Ԁ� �#<k""z���Q��`�Y�[�`J��K������$��M�{^D7.�=���7����σ��p�i����$�^�b�^�n�~V���	��J���/�Mn]x����џ"��Z���l�6�4�e���ȞL�7(1��7xdP�.���^�Rx��#�n^��`�c���t>.��x�X����.�	ڇ�����J%�V�صaf̘�b��f�g'��_��~���E���B�,e��~���.X�
<�O���@=�F,�vU�6U����zy\$�����������w�t����ǖ�.Ah��F����F��IBt�E�U��S(�^Xca1rr��G�a����s;\g�k�Mg{���]��g��r0������AAA�/FV��t����:�{6|cy�Yg�vD�ۮ� ;�J*D��H
x-� (��%"����h(�啛H��q�&_��@W�i��OW� Th �@{WWS�Ƈ��xԵ��������cN�۫{��bW�ι~�≟�?C��,x���Iq
��Q����Qx��s���7���vvV�Av��)Lh�Ӿ���,s�N�&}N�[O���ϵ���� J�?�nO��_?#��R��-��'@��w��!�`J__t�&W{J��]hms$�i�73�i�3$hPxR���RH�nM�c�9�{eT'M+�pʜ�p�މ��(�q����$�����:ZGw�$��n�������:� !���b��V���t'���N�쁈ͽߣ1R:��rC�=�XA�#�s4 �*�`'>���.e�ὣ�ǁc!~�fs4�����f�Lu����jk�7]Sv�z�6 q��]`��׊�s �kckV�:�(Z1J�7`o%e���u�VE�/ N�I���]~~ٚ1&ܘ���R��^	����p��'��бy�ޅ+�m=Y��qZ3uH�5n������̶!x�B+z����g/4N��\��6�%���?�3��?�)^�F�|���g��ܭԇ���\J2�zУgn ��A��S3o�<�~g�I�j�rѮ������29+������uN�����AA�8��7fb��	ş?h�xyI��_0VM4�	`w�ZtvboS
�f��=�PS?���b�ǲ�hO���(��V�F���]����=1rs�ja�@��3,��3�ÎR;�I}��f6K.��p���F6g|W��<U�lei�1�v�

 ���)��ǆGm��mJ?іA�o�T0=m��z��n�S�le~gexoA'm^���+���@G��1�ɬi�������%�Ұ�ԾЂ��!JS{`��DJj0G͞�ʫ�A���Ol�K�43� �B���zMA4i�P<Tgx]h����:|	ޛ9`Wj<V�	e�_�g�	Wq0g�Y3�ث^�����6�UR�EG�O[��Ui���qn�K��nN"�?�5{�c�����u&�h̻�C���P����P����.��)2��������5�K��	��Wܩ0��d�.>ik3���3���X�s����RR���Hml466����Rp�hp�k�9����_TDeޙ��x̐�H�<bo�]����Xyӌ@%{��N�����߯��c=8��m����nA�Q�e���3�aQQ@3MM' ^�m��yW�<������g�+�������O�B���@*i������s�mAJ�뺻9;	�#�&#���F�� 2A�I�����D
��2���4�mc4梒9���٭�0��@����`Ɣ�<m��!�L�Xt<��Fuӽ�W5�]-�g��Gnǩ�p�%ee�������?�J��,�)�
�-Xv���.�3v�^�%�6���|}{�m��YC�%�ؿ�߸tzPb�u^��4&�=b��W<�4Xjo�xݙN�4RWo�':B%:��T9�k��W}}f�#���C:�-�w���9���*��4���&��2Ř��<���(��#���Ա+�X�!v9��A�'MVV�~MvvvYZ�%��A�Ĳ�2�q/�*=�@
�x�n��b`��ɘ�ک��g@9�C�v�T!p�J�bM���O��A%��4���T��Ay�����<1# M<nzt�Lc&Ki�v����@f(�j9��:c~��k����:�KI.��>�2oT�M�
�B��k�B)T�	Ϸ,�R�?��K���\/3�K!� k\��N��,?0����:�����R�PivH�������Ԍ���©��X���&��^6���r�N�N@�=*v�����>�ҐJ����,ٷ���R\���\'�xZ E�� ���2ٴ���;�,� ��OC�qosTTV��,M�S�׺X�2���(��)�6�ѳ�b�0�0���)�1vt����HT�r�
�Ja��J���]S�#��|�[�-�,���ز�D{�oǃ%���]�ݘ�9��-F�f`���TN�,M����pl�RNE�����ڬbe]~�;������^�Zص3zt쫮ڕϥs(\mj�d����H[]VV�1uY*���m�r�{{���ʸZ; �/������	���zuM�s�Q7�'�*1�4P��O���]����{]��\iD��&A�ë�.�������v�6�_|*=ب�X_�nf����Zu>lf|�|~�}�E��Jn��<��,]���^���� *<��fZS�7�0�`����h��_G� S�p����L������`>�%����3Vk4�
��z,~�	��2��e�])=�(�l�~����������p���g��m�e1j����<�ݏ��%�ւ`@�>v��%��ᥙЛ���cV��֍ˌ���ZR���QI~�t,��.�o�bm�a�҆�_�9�ۨ��\BՑ;}9ߍ+QK��[9�$���rt���������.�bo�-�jE����<�}$ω�l�(e�d|4�&��,/���� �v� ���-����G�%0(ʦ0�.0�̥���5L}�6�*�}����$Ad����:<<Ja����c�|�@��3�uG����R�X�>��v5A����W+~:���3>ۣ���ݭՍ~c�<��L��qig.����9�t���{o��� �cna4����|aa!��0ʙ����[dD�������2�h��)�P�iD�{������)���j)�2_u�Q��8�2_>�͈.	�. ����R]�-$i�R����<����DS}�{g�������i���;�N#hZʴ�@�<!������;�kƺMm��ۥ���DM���U��76�{�5t);���qB-�=��h"�����?*T�팕|�����%�ɭ��.F����Ι��8YF1՘K)X(;SrgN�����5E�Xl�֧B���S�ʌ&����p
��0��Q8���(�?���U\��
�������f�����,Z�U���l6�@�T �c���������%Zv�BDtb'hjh�����H�5��h�mԾcP���N�nnnBxMkl
�<�ڥұd�~�	���&���tE��R9���VM�J��u}ؿ�7��z�ee=�5lg������Dc�+C]^" �D�)^>�cdj)B��vn0��:Sh��J��q�Yr�����b�V;D/'�A%����#m�z� ����v�X�!F��#P.�/�6�`�f��%Hk�I��,0�+����'��lJ�Ţ��_��.X�{|о���%��l�T��(h�eØ�]��ʪO�+g&8B�:Pʠ�����	M���Ak�>��φ
�P��XeC��B�L"��?�U�v���i��{�~�Iz`��: �CˋJ����Y��LLEh�m4���](ґ0�@%k��m�HP����w�����U�����2(��e �<H'N'''��DI��@�L��yb����K��ݪ��>�3w$$s�&^������s&T��U��(��{����ba{�
�%�!�jk͙RϮ;�[B�Տ�2�*2Z/e/y')L��~�3U�C���h���Q�b�KMC�B��\l/ ��5c��-�(i(�����H_f!&A����(�6w�>H��](A3��O@��5{G��q\U����^b��2Tr���I�%Q|����R#F�7t4������i���[ǘ�>�髤%O�IW644�(oU�^�"pp�<�]�;�8D��O�6��T���4��B`�R�w#��ߌ�)� ^g͗ۙ!�Tr*'�u�fhPA��GQ�z�l�ڎ�z�]���ES%_S�9�=fՑ(T���x�������{jT2@�5���|Ҵ�&�������̀�d,�`���Շ��h�g��+<w��w�na��ø��g`�m�p�` I�0'"���ke|d�H�'�}_��(?q�H�{���c����o����B=��|3_T�	�YS�;>���{�c�܃,��* � ҍ6�}�5<:JQ18�z��7�n��GT�0D8=�e��f�bz+�b ~~�T`�����K6���6v6^\S#��B�A�F�<%���E!�'������A+Lj�762'UbB�c�{ �ED��$XR��l;�2@��T��ew�ɝX�1"Q�ͺ���5�cpz��P���*>[�]\�t`vl*U�<	��	'?�g�TL��~=��2%}=.y���F��M�Y��o׀��	>Y��G�|J�t�y
3A%?�=`u�%څ�7-�=	���Ku;1\_%��N�:6�c���3ī����*����\u�S��]����i$9	aW�J�+��bG�{YJ��1Q3�|���h
�n:9j��ȏ��Y��˶��=#�p����ե7����Č�2Q�Аl�1�X�B]�!U"8y������
q�}�ɔ毯Ӡ��p3=���y��K�?��&�7��V��ttS�Z�ė,��gW�F���xhU����L$�g瞯	OB�Ǖ4���H���g�}Qv�a/N��w\���n�WG:����|ßO��!2ɀFXhE�M�wF��*j���80K[�����
7�K��ă�4U�.��<�>��]!��8Og�=����o6�M��&�9�ѡ܄kв��'���Lx�:݊�2�-yNC���`| T<"�T��a.$�_��5
��p�Z�m���9&A��	��!�]Q�dt����ǕD|����o��Ԋ�w��p��������P�T��u��BSP8o& ����{U���_���xma�M�x��@w�Y�&#A����?l���b���n`��NA'�f��qzT[:��AS����"�l�0 ]Ȃ�(��6�訩��l9h�����-��9t��ɗ\��,n$@k�D����N��k�]���J�e/L�d2p�8��r�< �Ek6;1#pY�z�7��u�ɼ������dz�XI�0�4I�(���% \
â+�!�.����q��\��ta������-�M�����H���x�o�k��j�Č�0o}�O^b�ӊ6�6y��wCp����Ns #U���6��h��hk�����m��d��8u�mT׎.Y��uy4���J�7���.=FP}�	� K�l7�a�]�`_}�`n������G����/�/$P?WVh/��WdJpYYY���hW� ��bE(Zp�v���x�v7�/���d�IQ/��t3sEV�F��V��s�;��_� �Ub`�Hٲ��e���Vmv���?t[M/йT�ll4I1i�9���
 ���e�QUL#T��}�UlJJt)	�3�}�D��CCC!~���t�>��k���^�Z�!Y��ℓ�����D�^R�GH�2��#�6�ҩ��e��
��O'����ކNt1A�c�E(｝2cݯ]{�]M ��iT��ZRG�c�����Gn�����8D~z�
�,�(��f��4�}з�vȋ�@�gB��˛�О�qm=�������]�������>��l��5c���H�OwԸ�X���K�=�R�c4��"t=:��J�fJ�FY(|�;fa�>1�ժxbg��L�,��LN��C*K߃/�(M=���Bx����W� w��TT��7v�m���IJ_�H����{N�	��g�+�5uc�'cwW�}hll����?�`�� �<�$����
�*p�����@�`@�.%@w�puA ��Z����+
"΂&�8�x��$��oߓ�@Ntt4��d���
�����,��{S��P�%D%$�s�n,�1s�@�����v�9ڄ�����w��d� �a	mԶ��W!W�#۟�? �4'��>s�=�D/%�A�ľu�yÃ�/��V�Z�D�k��ݟ�ߒ�3�c�iq��ن�!�3؛���Ƨ�|9���(nB&dx�/��)��.����-��[������1�m �kp��ۓ�O�M7x�Ţq�d���!�b���lgRjw�dyz�-LO]J~k�����*�qt���l����e�ͩ�e�Ϻ�s�[疱�0X��>������!��$�O6~~gs����:''��arw��)��)�i��RYi�[+���� �Z��֏�e���&������&��н��ڜ��Uc��1�&��z�ͦ��T�v����-:\fC��ja;����)�?��G?I�`J���{KbO���ƨ�y'[���ϟύf�aR'��v)@ag�n}���)eHsi�z�?�Fĵ�`եc˗[@ܠ�`�&���GH�"`
Z�W�j�}�51�dՔ���s~���xT��@���^ccc���gz�Di��D1x�D�������P�2�+R[#]��wO'6��
66�?L�̪�.."-�#Ԩ��P����V�wH4���,o�+�+�87�g���eT�K�G�p_�6�8ҕ���f>��-�߁��Q		����8%��9�X�9dX���
������m�'�����18�7	:X�1'ĭP9��݉��p寏�ߩK
�Jb�(� �NK!,��S�Pc�h;��� �{#㣽��;�l K�@{��m@ 5������1���Xu�Kq�����I��@$t��"ܓ��T��[=��5���B�3����4K�]T<9�4Z`����b��p6�~���\��!�����>M�^~�p�Wp+���[�9T}'�鐘��V�:Ogg��$1E�����_����$A/,,T$?�Ƥ�j.��#T9�{�k�J�B��������)�51�h��YzzzA��$��u��)�C�z�S󄡓b��0+p&�*�ߡ��y��pA��'�=�$�����irF��$�������F�8����S�Ͼ�B����C���z<9���j�3�c��'@�r]�D�N������I	����t^ �r�
�x�WN_�!3�@����?e�I�?�S���-E/��H�$�ffg�diㅇ�-�	��ovM�۱���L�3�֖;���!���Ig�D"�b�]:��"*�s���w�z椳�����C ��e��(��%����	�<Y �Y��n��*���noog�;r/u��n�L k!B ���T��<�U|H��������/Q��V���H��-8F zGq./�7Q��8���9[3a����|��X�s��!����F7�Eԣ~|^k�z��CNΥ8J i>��&24�P�% 3g8�_���, i�Y�2B�K]XX(7l)�+/��K���D$9������f��k�o�U��U�:�/����X���-�w66�!%�=�%����XÜ�b,�̑S�<Ƚ ����d�q=�?�����>���0:��~�;y�g Jv*� ���(m��G7A�A��s�C�n]8����2���Rr�
��u`�y疍�7ҷtr�uy���|]Θ��=�Z7�(����O�:8���s�<��M��5z���fd�[ �v�8X�m�;̓��k�oXC�++Й{�ZG�A��pV�P�0 �Q��Lu(�������E:\�wn��� ;XxX8��Ӓ!�f�7W�X?��-���=P��A�(#_c��2w>B5^�+�����������>al�]C�����3k��^7Jp�o/]a�K�'�i[_;�3ޤ��i�pV����`V
�"ȼ�����$ψ��W���7ڄ��$d�w��lh-�p����U� ���zC����b�H%#�6��֓Eo�{
�9_>���G��d�8�u�^<�Z:�*���9/Dj�k}�ϓ�l�p��I��W�|��{�Z]E��A���7�"Ӵ{���0�P@�y�~<�~��'���I���B�T��Y��I�BNzg�@T���'S'��؏�{c��5�v��=���
���KN0�֏�2֗w�g��==%Zc�R��� `�����mü_x�L)ç�)&B��@���t!�,Ύ�]� �'�D� �vh�Ny�`��P�����b�9鿦 H�?�\5����U���kC�iL63�hɮ�C�hZ��v�i#v���[�o���4C ��-:�hm֍������L����^if�
�y����}}��,�č��}OY5v��K�]��8��	?!�������I���;6��ӡ�nM�C��C��Xʘ5�I(���T"�ǃ&�h(Y���ЛF��`)Rf2�[��Nb(��{����]o{[������6��Io♣	��{�醪��j�ͼt��r�+f6k`p��W^x�?�we-�[bޒ7�*jq�z��	P.��Ե�����̺h�L8���2��$���=�c�M5�5����&��=Y�<ŏWy�v:::�ۧ�a�H
;�_�t��ְ;�5׋&�L^�#��u�������8�B��>:�^1���^1/$$j\�y�|$�g������a U��a����}A��v�kB�-���[�_M�h.����&@P&�U��vvKf�ޝF�ϥ`�I����'U���M��csuv�� �-�:�J�e�ك����VZ����t+]�msM�ab�ua4���Am��|��������ʭK����H���x牝����P� ��m���[���<�8F��!��,E�:t�
X�mr	*܋�K��#�qA�#[s�̀8���ƝT_�����R���4�z���&�������3e���8�{�5�ݝ�=	��$I��z~k	�O�9ד⽻ɼ�� ��%��z'�)ICß0Z��*T*
?H���Ţ�5�����m�
�e�F-Z;���
�|ܺ��~gY�y28�����=�&vȉ�,&��� iŞ���?����b��|v�����-�S5fFC�rO�R����NS}EA�tjVf�999U��}nU"�U�@�$S����� �2�������$��r�[��41\{l"�� ���ߍ�G����Gb���]|�p=�m&N�����:�i�U>��GgA�Oa%)ƾ��Ԋ����pCZʂ��̘������A9�
e�$�!�<�����F��y�gy�����ű�]m]׭�)�|Y;�2A8 �^J�<t�zYjwt��ޛ#'��~��̭O����5���'Њ�;?h�Ԯ�l9Qǆv��y=�	���"G����k�r�M!���N\9{�������o}�����""M��;^�X�v�Gk^5�OVv���<K�
ͳ�����d��aG~aw���޼�<�3$;������bS(#�v9��N�2�C���t���D�6g�'�OX|9$G�����ucK��n7c�w[��	3S�ܹ��ֲ��8�n��'����D��<�{�)�����q5549K+v�M]�o.��8�D9�a�^����0[�`Ε��N&�ز;��I���|�E��[rCy��1[j<4�'1��O�E?>ܨ(�t�u���.j��Zw";z;�%�w2�¡^?�{MJJ�\[�2�t�|�2�;�x]�����q#���8S���@���Ob���g����`�v�Q�^�ݻ�QZ�0n�qU�z��\v��Z��Ib�ǿ����Ҿ��V����!y���	d�˘�Zƍ���jə�_�4�|��:��<�K����꧹����E�8�g�`"'���^pXXۗ//I���?g޸pD�5~�j'�&A"ę.9��ܨeLwc(0i9����R�����@s�!�6q�t�]a1����v��$�q1�Jy�n��+!��jv�nll4��Q�L�]�}���G�����EЪ=��W�s8��t�1��n�x��L�[}氦}����~���$?��
w2��M��$H���y���mN�10eR�dZ���e5:�q��H�<3s�ʊ�I��4{�gN4�\�IZ3��V�����	�y
����_Q��_���y�|*>��+�Rϒ��8*˷�A�(�4�@�Bv��j�E#Z�M�T�ё�I�#x�Q�|b	F�c;{6��o7>6���C������dܙN����ݍ���ťU隯���8�4���5���O���(6jgvb��-��M?~j�g`����D��Y>0z���۵��3+�oKJ4f:.���S���:�ו.��1�ʙIIJ�[v�0���(*��ٳÜ<<�

�dP���cA��rK����Aܴ�:����P.�;@�E~����Q�Z�����^MLqrq�M�������;W��!�.����Π&<���xT�m����'�������U��UFF��I���?��������s������� �9xy���7ͺ�s���8Ǖ��j��af�=����-�y]����ѵ'��b5c����i�}}sL�x3��(�w�^5rIb�vF}�c�� N��s�JJ���%�=8����{u*p
�>:��5�I�;�z����c�W�ط]}H��ϲ���QѪ{�����5�!��㲩~�( XF�8��^*F����C� ��O��>Mo��Š����"��' �2��@�S���"��#��#G.\{������%��0��p+h�M��%D�����ㄜ��?��j)��`�,f �j�h�B\l�}��(�K�@�YƓ���^0�B*F�e{�����XD9�La�w�(4KK����oԎ�$*e|�nS=�T�����U��d��#�a40��
��5�6۱c�ʛ�ę����.f��%��俣^;2�y���a�HtL�e l˛>JsѣT��nIt%xlY�n_�k;c�`¥�'@My�"ݬ�2�>�۷�}�\�S%�=�� ���� ?�G�m�!I�gg
j`�z���������Ź��	���ߗ�oKHT��n�@�R�02�$�gNM���ͻ$�j�)x��k���$O������SqO]Cc���Џ�O�aqP��G���IOWJ�BUh�\��_���^� 8�3 ���N���d��cH�Sȿ���`�z[�N���d�/�P8�^��\U-��q�����i�%)�B�1�u�C�`k8�����ۋ��8U� ��]^�vU3砊 p$---��� Q��W?,�\���I��b�c��w����\~�����q����\ߕ��{�`ii��r�L��yz���p��tt�k�gb�����P�y��'��{{>T�$��8�;���>��m��o�cÌ�^0�A���`?E����񎥕U�ׯ_��������8���S5ե�"s�`ϯ6Z������n�2���\d
����'����hz�J����뎧����hR�BF�&�3�약U�쑽IE��"�ad�Z�&ɸE��[v\�w�U}���?�ǽ�}�����:筓k���2��5��ܖ�!����pX y.�#��9�C��e�ےA��0��ڿ@n"��D���'Kq^�����=������֠Cl�M�E��>"^� ��k�e�l�~�?��G�J+)����Ġ�����?a9����.�`��'4*���nL�.�rQ	چö���NW|��8Kt�Wlq�ZvH$>�C����w$.k/���p��\}����@�ߥ[kkk_x_-<�}�D'c���ݧj&�?B�&2��B|�]��;>q�G"%RT�pH�Αe�8h����$�Б�K�YS L�%��c��N�H\�8�(��D�A,+,{�U*��Eq�P�5 �=r�_�D@�����#;��)�<�'��l�@�<�tu�؟g[��٬{����_Y{��s�akb���:�9�:,�E�mA��]9٧K�C�h
���p�d��눧PҮM:�,5��S�O�����{�D��S
�;�R�������(���JN�
_=�$�U�˒��,��^�0F"/�����w�	��2V�!�͐�BnǏo���}�H��gA���4��a{Կ�ƀ��VAw
M0s�Q��i����j�|��g�MJ�X=
G5 Cd;������y���6#­��ק�����{~A~�HM��q���) ���9`�3�U$|@dJJ��k�DgYbjQF���2]9�rt%����Pݽ|y:���������|��=b;00�harj�����wl���՚�����dsz�|p���ZX��tBGg'@�^��z /��s��F#�ߝ$��P���5~�ˣԚ��}^@jqQQS�Ug�fX���W*���6I�'O��U��G��E�3RL8�`&zl���-ܧ����rj�`������K��(pi���������@�rUU��O��$G������MQ�8��>a� �1jh�
:9z{
��v������E�K��B�>� J�(�zR����6��OǦ���
�6ϭ~�S��- ��JPd�;�ł�d��+'�j5!�$��;J��#��w�޷j{�����v5)))r�_������^�1�����r{�=̏������G������:��`�*Er"�[K��d���|h�-���ͺ��{GTu�Аcjj
�����Zg�A��_,���n�3�O%�w a��p�5^7��VB�F£X��]�-uY'aU��<I�OG����+��b����ሐo��[=���t��j���gV�O��&A$:�gKp1��'uk��R���8��^4�S@:��F\>���K�5z����Jl5��+\�ݖH�G��x�|煿�i���r��������qی&� Rƈ�#��'/��W��gg�������� oI��&�L���M[[������0?�����`|������n��h�k�.q�ݳ�Y,5���Db \�1�|r��:6�֨���FĽ{����n?qf
7ہ@'��=��lG�}}��5��[z=��jU��j"Eߩ�+$iA��Wu;��[�F�O��������� Ʉ���� ��_.���Յ��1Q��7����5�o��EԿ;��X���oLBP��E-�(��9'!�j�)C��8����'���>�V�3z�����!&9��h����μ�n�Ϸ�KW)��w	%�wp#�/�Nv�A��X���U�DE��-Cю�~�BX�T��L�2��q��)�ęKz+?�I#���ڧ3����+aI�#�ҩJ�	��`��8��4z_P���LB[R��C�ᦿx�YtW<�uJ�a�ˌUuIWq�U{|%%%�����&�25��|�zb*+o�zU�oc~:ʛ�$���I*�>������VVV~�\�e���#����δ&u�ٕ4c0QGE��^��� UUgzU���*�I�y!;�@w>\����ޯ�Q�o�g���[��GW._� ��$;���Iݫ^S�w?�j��N�9�����Y�����}kk����p x@����矟��?u��%�(�����������"���7�`|E9�賈#�S� c���cS�I��LPP�9aJKLL����p ��E]���*޿����e�-&ʐ�����ZlS��DQWE�D�k|��tm�Ŷ4bـ{(��kk�hik+��G#���n=F%p�!$"2����?�C���˅�Ę5�l���U༤�Ѹh�[�8v��9N0+���Û4��VV@65ejfL6E08��u�����/��a1���-LY��I�o����x8���(]%����)�&���`5�q��ʁ���ڀ��~F��b̍��Q�_��=W�O��;\/�j�w�e!�K��Y{*>:G ���^�1%��ISx|����M�$���ͨ�g�����4��Z��[����h6M��P���. >�֫J�t
A����ʪl� m���[+�<�����%D�?}�9�Ą[h���AAEM�(�$��dvY��i����ׯ_�S���5Il*�t��͹=�M ����ƺ�^�� E]��M����JKu�VF��ܗ��G<�<��,#�[�R{��+�23�w��98���ގ���FQ�5;Vk������wf�a�}����F��D�&���_N�3]��7�嗯^��D��dc��<���0qǾJ�b��f�n����`�f$X`�wц���O>sJ�b���6���"�۟XE_	z���������W r���� �~=�ݾ������@������\��Sa+�Pr�ZV��]��ff0�'� ��S!q�'GxP��߿�yo�O��\�@�������,�IO��aT���&�����;ҽf��䊊��U��~��7\f��k���A�B^����^^^��5�U.���=#�oU�=]ZZ*����������2}�#Sa�{*�l@����V0,k��Jp����3bsuueV�IF���88��9t�?ozAʂX�����d���vzn#N�n�!�V�E�s%}���<%�!�]�Z_�Df__��c��4,Q�9�hü��/ڰwp`��ӣ��/d?���h����G D,@4��O�¡/産p�w���(X��1�gr\l-������G�
�JJml�o���G��y�o��}� ��|�����]�P���w�^ި�3���ґ�d�@��aG[x�w�rϳ,Qهo.�b\{�3��Sc����a������
]X3�E������| ����)���A�fve��^��]��6��.�N��C�O�sOP����,K<�݌Z�j��-uCCÖ�kvvv��Lk�j~J+YY����%WE]����6gF��j��s���j������ȋɃ�fkkk��[ۊ��s�;�a���u|}���i�hʺ;���;	u��|}����I���Yj��x��� -��`I�>�[��_(d��#�܏�{rYJ���A����}��U�r��ے�B��.a|V�߼y����P�0�}x�r�-z�]�cff����n^�9*Ay���4�3���n����"q��j#�Nr��~ʩYEh��-�.�ĸ��k��>���'a滳�7L��w'���U���-9 km>;���}�3��CK\���r�e����gff.�l�+W�o|x�Op��u,�ĉ( �sss�⧝���xH��4�x�_����4t���bm�<���������&y���$����BFN�l!�N�_�S��=�f�FA�58Q|VS�9�/S-ɘ�W�y���\ni�?p�Y��h����M�~�����6_U`/������E��L��$���ۛ�� ��vÊ���iЮ����h�u�c嶸��B�4�����������h���g���`9I��1����9mYP��X/���g��S�bkE�@g������ώWk�%,<��4�@Gĥ��I���/�v�����+��{z�/��z�*A@ �ܟs���wog}*�"9bg}f����/X�Ãi�X�?/]NR��UG4��H�ֿ���v�/����qN�g =w�2̇�]JQ��@�����"qj�>oO�	�
Jʎ���y�==�Ň��edNzYi�����rpqŔ����<X�24����:��晘p���ۿh���^����v��#Ѥ��$ͺ5�� 0;�U�ނe��V�j��o��ϟ�+�7���]�������f�X�����#���[í��l|�=000�1=@-�L��Bǂ.��������	�d��S u�˘�γ�͋�=��R�==��ū��aTb��>�pm
ÿ|���: ����ݰ�Жdqo�h����7
�¢�R�����������Qw�fF��� �,9�J7�]]]�`��<h��Y�Z���G&_V�$'�{w�"�$��l�w��<x�7ez�vE�ވ��[�d��yˢo�*��y��iݗ��XA�x���l��[	�����aA{� �xϙ�
5�o���?����̅�u����u����� �fxhk���%҈��P[��wUU�3~Ȃ����.�ЍD~���<>$N)*��Rq���Q���?���l__k�/5����oox��:d_
�Pp�~�nK���������u�G"�ln4�;
O��VP5���<U�]�J�����ܻ�{�Z��' ����t 3d��ǌ����� �����]]�j��}
K�D%d�u�y���5/:DQI�Xb���qDo���.^�䧺}c[G�<L�ؕO�!t�<c�$X��������P#��2mo��s s�|��0�j��4���L���r������H��"4b�/YQvx�u~��{��]��*�}��%��&���$�ߟ/�n���Epn)� ��&��ث蘘�D�MZ*���
w�5o"��@�ټ��k����{�p�9�30��mO��
I��3/鏜�ÿ	����E�~�q�V�Ѷ�k�z�+C�\���)U�Y��TN(n$#=]�`C�kC�m�Et�9�����C���/�`u�u�g��Q�m��>��|]Ff2�{90�,A{���:^�(�b��#(�W_(��D�[�_���#��_Ҿ���ڪ����'夕t�2qp����8!���<q�e��S@t��,b�-.��>�t��(�J����%8��ٺ	#{;(�~�N,"Pr'J�zl���Sl�w���j����+��pB�����յI�����S����ϥ*�闥>L��7���=I��|KA�d*�C)::�ӻz��e;��B?�+FЕ�r �o��������*�
4|���#7%63����2�{�M����ܗ��vT�%�|4,ހY6��� F8՗�YK&�*���h��}�X} !�x�eL�� h�0�����4�|-P����[�m�ն��B�rIm#��]U���aB���r��8�	����p�_ �}�ǧ�q���7�)����������&zX���(��}E���ߝ�q�͑L|p��Y+ՃE)���(g'�xؚ�v���L��p�Y`�Y����[�ٹp�WIQq>e*i���K\��!.�6�b*���~�%�O����s,b�n^�w�[���m��P�{$��l��C=�*Z0P`�h<��5�(�[�����Ϸ�\
Ǳ/�9tr~�f­ۅ�\�AK��f��7�����m���x�>& Bܻ'exh�AZ-$qA6ت��������D��fK$�R�f�f�j���Y+��2�-#U�~j ܰ�d� M}�V
���wQ�,�q��cJx3SLK�b� ��%����w�1QO���~�����7 Ȫ҄ǰ8R�А裒�Q��
6�j�]�����u.6�&Xޣ� ��hS ��i�����Go��}�ݸ�	���2�z�O�ø��&w��Lݍ(�#w4�oď0Єafg?f�+**B_��%��Vڈa�IF�0���5p�j�1 `r��*J\z�j��:�}�0|*�^`ι�����Ji�e��vU�kk}���I��hގh�T�{{>v��I�)e�i�f R�ι���JHpj���Z�?�!_0*'��W�k>�b�8�$���B>��D��:��Dpna���ehf�a�k\�DI�շ���#�3�L��@��U��ϿdD���B0E��_i2���?��1|�=4,d�(�}H�rr�����F��'��#пw�8�U3�#)===��*�� �)��M��&�jgee!v7�Ɲ�'�?>?;����&v䴆���5	����J,)��%�UUe,**Z���RN۪$����۱y�M	�V%�X dQ����Kީ˻-eBW.�C�_�8H��G���/lj��k�ΝKߞ[Z�����Y�<t֤ݰ�����{|<@k��lR��wr�{%�vo�Ȫ7��Ǳ�ϲyUA��p�X+�����[�7�����G�O��pm`�E`"�� p���y3�n]8�ҩ�6`����r�M�<���~�[.rF���x[Mv��v����Wy�k䋻-�]���c��[��tl9�е�72�K�oPvC O�5�����9a��)g�Ţ�RŰ|���[�fj�r������\Zz��"	�KNî�� �/�=��`�!���AA\�����PM��h�g%�O�XJ�}�G���&��P��O��>(?�����MY�QbC?�wꬹ�:���D��Ǖ��&�'���8�8���[@Q�z��6&�M35+Kq~a�8�����α������YĴ� Н6f�RPPD��2NLL\���1}��U�����_&V-���T��c���-��;�������D�u#Ew���mUUU�Z<5{(�<-��ee�k�2����k�! �l��Z�ybȘ;�4 ������!�h����Gv��HJJ8�(! 00���@t[-�Xu2�D�5nwm�DSE�&M,�:�R��U������`���`\�����ֵ�2���1b�i`>�yp	���^���Kh�~�_|ՠ�4�V��1���c�M��o��m�i~ɬغ�48%T�`�#��P��a��(��E{�?�@���Z9E�X!2�s*Fwn4�Ʋ�f���"��|�F�'Qٰ}fff����v>Z�q�[�4&�pof�4��wС��������fI�~s[[i�!�}s.o�������Ӹ��@T����}=˵�c�Z+~'77� ��斾�J�9��H���<�\*)iq���������9���q*�+�KO@T(l^��s�^D��z�ܙ�aAql����.��	����(�5x�BJ�/�{�*�Om��N?P
�*��j����oGo/��K�Z���e---=Q�	0��b���7ֆ��TD�`!y��ď.A�	��/%Hf������8T��M�H�w1�P�^I-,Ԭ���Ӳ�k��������F�)�܇�;��RSS�˕�H!⹖곞0��vփ�&Mطdq���S+���r��BL|8����{z�'������MCe�ś$Ǐ��m����:�/`�T�4��:�-�l��%��7�p�j\b�x�-�.J���',@�	��:t���mRD8�R�!q���U⨲�V����yK�E�R��GX���T��I�x���+�Z8�~O�a����2������dld����t����A�n�9���R�a�ý�Ü{Y����ݽC�M<n�#�?��O?����#��(��5�W6e��}��`ێھ�mM�)��"��,����ޯ!Tś�g����l�n�����IZ�r3�z�e �b��b��/a���Qm��A������f��
�f�G��Pu��P��r*+�X�'"p*�;Y�Y���2猩�|����ᄗ?Nn�u"�T�R����u��^���V�Tx�~v��w=-��/c=������TL��]=W.�t�yv{�0e_Y�
1�X��k	������1��pa~>��E���D�{�:��P���O�(sL�f��ê��~��҅��n��?�a��ܹ3@�|I�ߺ=�ZW�������&&��53ӏ��
K*8=�Yiwq�t%����.}����\��z����z���44j݀j��YR�|7A�KΕӏ|>�Ӵ:�ӣ�xq;zhb�݆��G�"�e%"��N����+@����+i�v�,��ᱦ~��Wؼ��b9ϝmI��=��B �Z9�F}�6A�5q�ړǙ���X��JGun�],�leP3�v��~4���(��
���D��-fy�1Ub\��m$9,��=�
d��h1��Ǐ���t�'�%�֝��c��_��73k�9�S �EG����ʩܝ�N�)��es�O��7����5<S3�������+Sy�+Z&B ��Ž�{�.r���/��mi��`�C�#7�'�[����=^0Ү����d��]n���otv6G�?ɂ����<L<�U�;�#
g1��N}G!ُ-K�B���G�Y��o#5�5G���t��CUL��4����}��������C>�I9dK �57��5�Z��MY���M�m�0���$�Ӝ�l�ⓐ��?�Ȧ������������ŋS;��Z�3ȅ�]�ݲ����1��圃��;_������j�΂=�44Ȃ0���0%�?<n�5/ +����]櫬��D�
!!��w��]ᯁ;�D�$�T2�U��i|~ݲcyZZZ�Q�JMsgf��,�4��<����PH)'���E'�O�G@��������j�����e��'z D����������ջ��0{lv�N}���h^W�����j��N�ƉG���[<c�J�}mUj�L;cl�èP�?�U��������2���¢�6&&��ؑ鶔�T$�g���#U�i��jP�� ���U�jW:,[+����by��/��������?��߲�hM�  "�,A��C�c�˞ �v�]]/������.��:2V����F�~�����]�.�jim�JUspX1�����l��!k�Y�E�P|/���<׿q-dhܠ�1ݟ�En���&v�S8��:=���ã�kL�l9��&����"ʹ�&��������+-�p���c.��ݻ�1a�����c�<'#�&�F���HƂ�q���	ďX�*'�t��D;w�x��>8�EC���@�յ���n+
�o9�';]��\����-gѠ�B�d�8�INཀ3#�*��/Iu�J8��	O�'f"Dr΢iE��t��ZS	�q�	�/e�Ռv%�ʅ^��_#y�d��aUG��í�=�`�x�C0��=�5���K���R���#'��@ Fw��n�2`z���ᄵ�I�ǔ�����2��J�&���gp�%8LLL,��}�����˒~�o���i׊_9��\����<5�Q���2 ��W�7f۳�n�&0���]�`j�|vYy����6�k�5-�_C�EZiio�/Y+�L�����1G��/�4^�Q���uTh�oa����3�%� 	D|w���w޸��R���q�Ƽx��Q�e�1`E�?����AO����`C[�"�z^�H�'pJOnAj�4x��	Pj�5<�wG�-��di��D�����p��!;ާ䬀�,GOѾ1�T�|���#i�22�������,���a;��* �a�G.�F���/����b�G^�����mj�y� ���htߗ_"U��jv���@CE�_\�-�?d_���㴻a�����V�۲"&  �b�6t���t��c�o`	���K+��ZϽ�,w͖�p�|S�~�#ט	p�$��"GШ*�y�3�zK�v���>�|�ᔀw��Y\��#�N^\�"�`���h� �΢�n�=+��$�2F-���>O�����ae�-A?A?5e帑�@���U&w�|�9/�����*D\�uy�ɋ�Z_C��ޘ�fEKW�#[@8���%R{�����[�5�!�C����A~a!?�J�����v�pB�޾o�H$���aZ�����K�z����-�}�����ŕ�-5]�7&��� �rk��(���
!������y�=��*�p��S��;2G�4�+u�W*P����z;�/����b��S���i1x���`��[�W���4i���� �m�]���N��ᩫuwsЎ�\�+v�Cʶ��#���z���Ǐ�T�UTn��}ق~���S�q�'�IH݆�Rjړ].��3�.��'Z��"��y���z�9W��bR7�j�j���<�|W�;^����@?b�*�FO���)oe9��7M�������4�e>gٔ�~�������UN�]����\`�N,c��!`���5 �=��)�M��!b!�����25a�B�wLtt�W!��C���KO�g�9W�˩n�~/���ή���?~�fl�$���w�`���w��@QsQ9,�n�2Z������bϳ�:�Ȑ��˰?�IDEE�1���4�����)M ���#m�ݎX���G�DD\��jI�i�	���i����i9^�Rg�_&'g�����T4�~NTL�z��v�i[@�,��]�6�T�E��(_�M��O0Sc9��m���4�z�1gl�_)�&԰�O���A ��l��@�-|�=2+���W�x�AG-��^�2ᖮt��C��i�$�t����Ǚ��j̫PLc�f��/d?X�-� gwٯ�m��5T����2�CJ��4�d]r뛚T?�(����&q��tX�?�.�1k[�,���9ⅿWp�L�ζ�C�E.|�>�|�P��v���~��X�0��^�v��s0|��Da��YK��o433��>���Vh�)��{�ǖ��2�;�0G%�#�*�L�Ό�=a��(����ٳq��@��o�9)Н���+ʏ띥�����;���� 7�4���~b�#�+>���/w�����w��-/�ed4vрTw[��&��-���W߾�
�ȁRA��
Y��H�Dqhq(�ź�2�u%�8��PRy'	� 4a�̛��v}X0?s��/7��hK��h�r!DQ��J#�r8�Uܾ��mv�}��9_ Ж^$}��*	.a�{�p��}�I�[�;��d{��)8ʑ�63����L�2?�w?���ʪ �$��N�����|=���o\�1������
�$R4꺰p\G��T%5�y�[(�ݣ�s��f����#%$l�]ǝ�[tB��\-������S��+?~��J�����j���b-�zc�Ǆ���g���WHFz����}Qg���1H�~*At����-����
�Y��ő����gT���$�+*�H��í��gՖ5�"�@K�������t��,�uO�>��Tr�} �Uv�@�������[���SY"�<�Q*���?�0�<������=|�AzwhÃ�� ���Mpc2�`.�%,�D^b��(�1�;��f+��N��=4~���~�q�x�^ 'M$�����l�~��$�hS|�I��?�ۻ�
)Ͷ5o�G�[ ���7B���1�2񫑜�%&&n{��s�j�uã�'�p�5q�Y&+OOO(g��i$|���Jsst�Q�M�aD/�G=�9���X�������q���g�
-m��`��Y�Ȗ�컛��� ��S�Y0��}8K�����KŇ@f����o��q++��~�>�$,��G��½������Km�m0):��Hh�t0-�+S
4R����?ďq����Pj�0���fVj��@)%������+���x���&I��$'�.�>�舸t����$��cJX��O��������IE��~��@���w?Mvvv�0'��ߍ�� �-�8�2 %%��e�X�.Ò_�Q �b�{i4H�����Ñ�is�Z�ɽ�sN�W՟&��O��w �O�>��Bz��d_��Uw_�]�{��o?啔^���Z��w�����cɞ�:yFV�<~5�4�{�v�%��j@¼��E���h���.+������]�%v�����;
����3\�w�%��  ����J�m��C��Ǻ�l�Ӄ%Cn�(���t'��S�4Q�����!N��m����I��<��;��̓`#^�fFtwgY����9D֑Rd����ݢ����;���a�>�%����N������5���YGo?i:(xiI���;�`���:����.曛��u(��-��A�BR� e}v0�Ȉ�s��@Oͭ��vf���U6ᆠ`��;�R����U&�*=;�"�e���>�9'?8���_;Q.wW�KJ���K����߭G�nk�V�9������V���2.Qs���ҝZ�yyw���*�:�iG�Դ�;~�	�qDM��D���흥�s��BniKn�;=}��V(�$wcm�ݏ{��u��?�����l��5����������G:���5�M�_��#9yǃ`E���;&N���ɂ,LV�4���`d;d�p�FxGx��{o�/�;��"-��f=0�{	��m���l��f��h�<�����fe;��t-$yf��!n�utt0��kV��ONM��8����(E��V6�H֨'x>?��-�����	*'�?(�1��e133��	�~���?�r�Mi{�]�������y����I�r<���p6:ߜ91�DĬ�Jru�2�����b#��R^��������tǤ�~y��02�lhhH/}�����Uʈ�D�;�>W57g:�}\@B������`<��n��t����am�x�fQ0NŞ���x�Ɇ.�Ǎ�8�yl�������nͿ{|�1�6�6�}*׿��a���t#��2����ަ����ˬdO6�x���G���d��1��2�\*2�;���6��s�5T�?�gٲN/yK�L�\}r
w�4@O��:����ln�����3&ם۾4���G��`zi���1b�jI?��a�(W�w�gdf���1&��[w��Dk?U�X/�~�{O*���IEL:��K�qwa£[1�8�����!9cN�_�Hso	:G��)8559��M�V����!����m�ۉ��O-��D[XXPaǓFWb_�<��� GkF��r��v�֦x���~�Fw��R5Kh�`��O$��f �����n��.���ROo�XV���ڎ�ҡ`�~��'��:�b�ڀ�PZ��lll���3^��]����^x'��=s�E X���n���Jʎ�7s��h����\-.���'��� R�?�e�c����)�ekG2��D"�z��� ��5��B�7L��Z�u$J�w<�|T�{p��9����Ԙν��12����Q�0ʪ3=n�vG9�຀�$A�ҏw�p�"a$����Kr�=�*'.�p��%+��iS�~a�J<A�
����~��k�4��͂r�+z��GW���� ��n޴e�Y�h)�\�]>�,5/�U^�WX#[�I���Ku0l�U?��7��D�p�"ݾ;K��IK�A��O���|dCI!m$c����k	�{�@3�{q��9�)�W�|hV~P�6�f���<�xL�3�'�|eQfV_C�Mè��_XA��2ׇҍ�ԩ��ϚI�QRR�Nڅ�ǁ��>�,��[͢dC9W�ؿ�������\�q����<��o�P� 5fu�X+�NT��M c��m;�ܙ������ײ���+ B����\T����AAx�A��������u*,,4�Y�#o�Xm�B2��/����E� q�71�Բ���b�����_�Y��qD�{�t�\�������?ԕ{�xJ��BA8�����u��9	l&i����!x������π��)fP^��f�R�g�݆�MƊ�ʛ���I__S@9g������f��<|�����i���\M�WZ�d�p4��d���G�zTa~��mKv�0��J��f�$w)n[�b'�IEU���'��R{;S�+� $�V�-E�cK�5���o�]����L�F� ���=���fwVU��9�9�;�`�Wr#P�Jn�}�a@2u�M3�����t����{P�-,P,R{|O�Zh��)�,\*���.���x��_7�J�MM/@_&%�K�ld���2#G-�>�O���S������F��̈8p�
;��m+��r$����U���F02I�d�'m/��<��tQLk+r
Kլ�%  �-9%�i�ǣk7��]��*_�M�)]G!/���7g��Ns��w���b��Ktadb[�sU�ocDt�ʪ�-�ۣ�K�X��� �i���~=���IP`�����au����������.,���I�������ذ��~ �B�I�$wA�� �X6���X��@��J��	ȗ;�u�\\*͢R��ƈ埾:z�+77R��l�9�8^ ���Y����3����Z���U��#p���y�(O�W��pywL^sS������َTe6DȄ�(��?2���u����^~�˗��+5��KlG���K�fHK�l(��ɡ0 b���w�	���Z�s�0�,���kɠ�RR�
073�~��gۙδ~�Hœ	#:�1X[f���ݕ��k�XA0�����W,	��F���6������V�ےŏ���S��à�]�F��_������Q>;N�YqK���z �~Hww�'�����9���p|\L�ij����<D�~6"J(?��~���a���R>�E�v~(��X!2&���;�5�����7#�ϟ_��J-��S��Gv=v����Din��hF�ь���������(���s�
o����CF]�(�������J�,�b�]e�������f���k<z{Jzے�%9GB@@��ynnv�q��;�~?��Pd��\@Ӊ'�v�3b�?���!������7�}�>�Dó(տ��4����Z98U�v>���9"�z��:�._�x��	�˥3��LN6u�)� �?�-4�v#��?���
n��6��[�H��9��7�V�,/�}�=#�S<K�V�%���z���uƓ�d۟?��9J�!��;�qc˶ʎD�x�D��j��nj����v�R��l�"������� l�S��� J�,�|i�D�a)�)vxQjj��z�L���h�M��/�oc'�'���V*�)��� 3�]ϸ+ӂ�AWW�<bz����w�.�k�tN�I�*�����/m����\]�l���^�0���|?��Q�f"lL,6��d����e\oSPQ��m:�5��¯Z���G
.�jPts+1�K3@�17��am�����M�@<
�_d�i�V�WR�!�<��6ٛ���>
w�jkΞ=+����r�*r�4C^�Vb78	�����B�1��_��:O
JJ�r��90��bnMݺ���X�;
6�~���ݮW���m���V�^d���Fs�!�D�Ę3z;9i���bk>������ �>�7YÏǗ>�8���8���_�=pqu�j�("�u �$�;ccb�����Mں�i��fJ-�hrS^ɤ:,��N�����C�H%0�Ԫ*�����m�RC>>>���U r���}%�*���!͛���^�~��־{��I��5�wy�e{����N��	|11l'�!$�dc�[���	K���Ez*�4.����������N���E�g��3���5&�n��e{k�5�+���������g���ə(
ތ#V&9�.|��{�z�Q<%.!�9t,��#5����1K.������%��K�lg:�|i~v*a.�����]=�^8��D�sq ����d����_Џ(".?,O��U L��Rq�����U1��r.�`;| ��85��Г���RbW��y$4���`�u湦��
<��<�ڝllbB�~�=jj�{�JS�ˬ,v�ۉ�W��u{�r���̯f���͢�޾�""lHs,��L�X��z}��l��ily[xp�9��� _���ix�	�����u��ں'�R�'�l0�.>�@�[�8������u��J ����&����b]-�&$����Ϗ��d�EVQ{`�f����UUU��+� ����Ŋ(�5��$�|#�ކ���.*�����05��U�@�>�� &�5�f5�~�h:\��Z��@)�-,,���鍌�gE�W�稶�[��d.᤻�1�ǖ9���m|���m��L�YVV�d�o׫�*.X{��ftB��C-�_{#ef��҃�.����>ne	o���R,�O���Oɫ��a�k�ͻ��{��
;J)�x��~m������V�d4��J�]҉y�C������ǍQU���vv���9����ȑh|���o(/�{w��ׯ���b���O�P�	mA$m>���~dG��
deb_S�G�|!=�L, ,l�u����cXF� �t�b���vI��g�P�Z��L�@��[�`z��#4�8���Qd�����c))�Kᬬ艝���X��A<��İ7+шyj�9e�y�<{������,bH>W�����x3�ATZ��	�>��(�G��V�ȥ/W�r�µ"`��.tG�ټ��_*�4D634O�bUv�o�r�#�y`E��js}>Q�,�3򌢴��;�g�ׁj��q^Tx����V���܇������ss�f�g�Oݕ������!�Wy�G_��͟6�ha�4�"''S{ni
\��A}zY^����ch(q��v�8pNɛ[�xfv���+��0����5r��0޻u�����T��Ç��D�_J�W{"O0^dFKONޘ�2,i�Gf�f�Va� p�!��CY�������s"q����.�������T#����AsD(�ȫ��	�{��h1����>o��D����ܢg���Tkz^��R+���*��-����L���"@a�J��j�wz3/���8�|��2�)��ԉ|6O�:=����`&ɝy��\��O�~������ˆ�K!+]S�5Ѳqp�r��_�����Wܑe�3��%�J��`�+_�>˴0K9t�M�7��@q�ѝ�S����$��,\�[L�U�U��#��(��Ͳ�_�%k���+���ю��������œ_���OΊ��߀���#2�����Zq������ ��K	�n*�<J����4�����1*���+ "&����޸N���������z'-�i��H��9�	w��
�|{"w������F��]���z=CC9L3>[���K�K�]����G�'[[g!��XY埿�`���b�XrT����
C%�pK��E*�ޏ�H�klck���Ѹh�_A�������_i֜מ.�P|f����r�1,��urvrB�u�ɢx�L9Q�S�o�7���/$꒢"^ݩyv�Z����U	cU�۸n��.*�/XY[w ]���
ff��0d��Q@A>�-Y��8���.���]�e�R�mǶ���HR����A>7�;�.xn��&M��ïƫ+�����]x�ssF����	�9�l��\��Ē��@��<���=��j�m�;>��Z*�<�V����1o�ma�qU�G��A�8��
@ml��/��/}Ԋ�Gvuu]i&�ÛF ����5�f]��G:D�WPpw�BV�_���?R�2�5{��-6ORz�$���F��[��}��ol�n� �`��J�[~@k��$i�̼��2�z�2�ee�|�M}�Vl��c�͵�`8M�~}���W�G�:��ML��p���j�C*�����	�z�bm#p��}��2^ c�|����C�@�.�3��ʚ���w��Ag1�՜�-�7��:_��D�Ċ���q�J���L� \�q�d�| �F�ttt�{k���-`���[1���47��D�kÕ�%�0r���D����7� �7R�8���)J�����'Z�*�z�� �n ^�������:ݫK\�6=W���� ���P�{����ĺM�6�s���������
	�(.$$���6�G�-��n�>0��.�e�@��F ��0�p��U���hq�2�1 ��7@{//A`Vxir�c=�����LS�87��B3ZN��x��ϵۜp]�T���2hV�9:��((�(�$wrr*���X��� v��pM�������k ����֖u�`g=��
3�g�ֵ�L]u\��^�AAA����hP�I���C�AJ�F�K$w		�]\��3������������s��<gΜ���"��#O �FYCc��a����
� ��ǜe2��̪^��r����SQ�PQТ	��Ɠz���}�b��Z�����K��¾��_ uwtH�ެ�Ϟ��]W��e�g?���$2�z�	D� i�zcjf���_�ge�tH8�J�����V��X���uᮛ99�~*R\BBo��Q����g�2��:m�E�ә봟�`�y&�FPP�T��;8���%!�=OB`��������2��4�tZ�x���������Z;D9)Zj�z3�H0����[]|1��b`��DT��[fVD�7� }b�����ua�U�9*k`z-}>4)))�W&Rƅ��]�WFb���ؔ��ڀ��\�)�Ӭ�����7�6L$�w�LL~.�����_ Z�=���5)I��ԅ1����*�UO�c��t�"�2qbmY��߳�Q�2H��;
�.��e�������n+c����9b�m�%��xݳ��]��=�'4��s�E�l>�k��:��/_�li�� �H/ 0��)?<�X���Ý�o�q���F��Dt�rV(���V0q$���U���D�_ʧOuO��6P''. HǍ�؎� �u9��;����)E�e�D*k�
P��9Rqi��2���k5�G�����m���zb��
�,`�ab�9��$����p<��4B��B�o͊	g22���=ns�8���ǋ�5\���R陘Ĕs�3ؗ��.��jF8D\#k^�m�^�'t>x�^��p�?��m/R�n`�.y�}�CT2�<,�����0�
�D�3���7��T^�JJ��{%o^�E��%�5����$o$�x��:m#�qT��?��
�uD���`
h�ސ����Z[�*0�>_���8%�x��Ӥ	�o#�.���l��Ug�z�����M�a��z�����i�x�C�Х���v�*��p5���U��O�/ �����hEj"ۖ-A@.Q(���ξ�\�����n��މ�������/���*�E����\֒������&*g�Vy�0�	`�@����7�ѣx�ٸ���D�Eս����dȳd�+�����N�~W<��v������ �@#� ��_�)���nz�TB������:J��h�z�Yj�P���x����<����1<2����s��Ya���	�Zf�i*�;y\�	�2���#�[�K��yy2���tŬ�?������	@S�edd܂22��R����"���@��R_��q#�&ב��]�L��\��t�E���N�v��,(�}|�U;��T=1�Y`+���k��eQUU��z�˚�)��SP:{�rݴU{)�.aoр^`N&	���X�
TF�7x�(��i<��M�Q�t��.^j>�{\\J5�)�,�.��܉k���)L�RDVnE��2����������ILְa)P�@5��ի�JJ]�Ѱ���K��y��)�NEI�P�
v�X���Ս����"x(o|����ۿ���@fƔ�ݼyv4)H�%�}�G�3 �-���s����"�ƈ}�6'ye��(� ���W�q��ڵT/��1�n���Է�x�]�p��.�03���q-�M����tv{l��Kx��Ve� ���s�.&�<�$}_ɒ֭ց�vK
����Ax���i�w�d�ۗ����qr-��1N@Ϻ�wt�ٶnӭ�#��̜��yIL
�fѵ�S�{y� �w���������ng,_H\����ցN(��$D�9��'���c�;]3��;�F����9o^���4�����\Cj-&*
7@������F�[O� ̀%�;.���tƑ�;u� ��NHfg�������X`����g.�z�V쥭3B|YY�̓��Z��o=�Vh���t��V>�.ئ��րfX���EᎥe� ��勬Z?���X��܃�8>{��/��^ZZ{}ZR��ó�~ojm>Tl��]	.6U�C�T׭1�/3����zb�*kk�p䩓'��,q�D����� �(��� ׁu1�����g��Ŝs����F���.����q�w�`�X���^��=��ϵ�k#M�@I����������2�/����lf?��6���hxZ������]���.e���q��Y�-hw���x����4�fq�d#�T�\����SD��e	�Y�|�07ϳ����v��%��.t0�h��
SǕ�m�[+zT����c�=wX��XmMG�<']�L�L.�,��w:���j�[||[��4y;�Z �C��9@�1�Q@@�O����!}?h�p���c�*`�b�Z<�ߣ�J�ݱ���[YԦ�(J����e����q��4l��� ��t�c���?� �rp�����}'b��h5�	&ڬfK�4/<������7�M�g��|��.`q��̜(��QvyN��yǛ�b�z|�7B 9�)�6qʉN{����%Z ��-���?�к�;�d�z��jC���H_?5�6�r�c'�:��n�%%%��翡��Q`<��1��M0�R�h�lt��cr�Lw�~n�����P�����R�J��h_s%-�� �*�z�����*J#ͫ ...�J�f� �WIE����:UjpDB ������26�;����(��s��O�a�(�ˬ7U
n��Ol�zO�Z��8c����J�����a�@�`n.��6R�"!	+��n�-�Z���O`����55��(�� ��Q�����e)�M��Á�6 �����C*2n;>�������A_Cw��8�s��GR,�� ~6���ڂ��,��ޯr�p���;���"3$��b��h4���\i��_'aŀ*lU�"�k�>��@�Tro�~�\C���P�m֜)����@�qݮ� a���^BtL2��ht8�>rw��a7�gl�3���O%$B��ƣ�ѧ@֒QPPr�F���2��-�����-�n�X8����
 ��,�d?����~�;��i�_������\����a��i�,�+�x\Ix�ry���t�Ƶ2��S*�H���;?�r�����P��ۗ�vl Kbae�ۜ=�w�.eE���8K�3�F�-���{��##e���`K*�0>�ߍ*����P�Ba8�^��W`|���'?|�;�0)�4m����"\#'�^Sd��PQ���d@�{ ��ba�J;��
�$�JJ��fh�
�g8y��݀�|���]ՠ�M�G]�zz)��;�2�>���U�a����:(�,�_������!�����1���@��R7�*���a9�]]Gq�����������,�!�~��e;w���r{{{����H�W���.QR������}����t������vvV�ޢ�,�i:����a�s�l�� ���2���V�ZN�u�H+r���Fئ���s��c�54L��m�n��-�SE�� o�8�8ͮ}�H >�מa���sq����Q���*�2��X%�F�Ӣr�����DY�@��t{���X�&��/�ʰ飤��r������4����(�7'�TR�����_7����ji�b�S�A4M��s�<~���
~0���\�m�
�X���_S��^�(l��зr����&�4��&�:3�iΞ�&e��=���¢zʛ��0���ǫ֞���y'�*�� Lj�H(�*��Uo��1? \5������W��Ne!@��7�kL�������$��m�w��c���W\�5���?X�.#��->�5\Eӈ�6%E�mӨ㿬�{�<�r�K+�'�[E�^�[s���'�+��1@PAc�C)Y8�~�Q���p��$��J�|.*�؀��wt
��4
���Ǯ�xV�摇@uh.v�^44�<�ڲ�|	]<ӡC_}����`>�T*;������a��E>y �z��݅�}��6V����c� ܷJ����<:6�n1C���׆�	6�n����vސ�%��ڤ��(�� �rl.����e���N��"�Q6�e���b?L�Zk�����6�6䨘���2�a
���N-��ұӘ���f1}��6TF����5ر#�ĠWN�g�
`���W`�m94!jT�+l�u���(��h�4����r�����>l���|Gzz��������sjR��[�Ɛ�O��풒��²^�YUoB�Rc�/ 8�)U��o3����B5�5��
�o��T "ݢ�f&qƔ�mooK�3� j��/��SK����L�3e��(��;��.8��V�a; �v+���?=�ak
����C� �ɫ�S�u��t�ǩ���e@�{wL�5�/"KeN�:� {慧��c� ��I<V戲��<����6+I�@{^y��Z܂���0Bu&CK�����0O8�7�W��W�����|�y�z�jk׭*Oh���,����*��p��&�O),��n����.)�d��ۭ��#��ia1`(�@�;]3~Ŝ�K��KBe���vO��z��de��zQ�0^Q��!���	QQ�D'�(	0?�����$�@5�=tS������MqLo̱}�PZ��)��f������ ���ꖵ���Ƕ�Ka�}j�R�:H�4�%}dɽ?uǀy;���mo�Mq׏������NR��ա�=7��|��
Bv���$��n��3W��r���w�%�߼�~�M�Wσ ���me��}�8&�#nY?��K~]S���a���x��)Y�ie^�Ww���ykXn��Ae��o��*��X�}t.�1���i��Ey<z��Z�R͎�B�U����Us ";@O�����̬,=++yg39�`2r�Zp#���]5Bdk�MR𱜜I���PB���Y���Y����1,/���QF�=��To���w�R�|�L��*��ʁ8ٻD�C����q�"9��ki0]�A �F7��l��Οn-��3u��Hk,`�EZV�~�W�1�<�ˋ6B�Y�I 1
(���g������Ц��t��R��;]Q��F������۴>��`��fD�@����CW��=Grd�9��6����t��]��� ��<j�&���.���)��U��H�ka��g�gc~�<��׃�I.P,4U��hz�@�^�[-l�ݛ��ǰt1.Y��`oG������j/N�[[ΡyC�T�'�8��vEI�+6�ί-wpv�w�jT��?�vB�x?X�w.�Q_���ׯ�C�`�+����zG�4���Yq`��&}Z��3��M��t�)r�0����3�P��_��O�N���ЪsDK�ڙ![h�0��g��d�eS�t�'�@��g�d��)*w���-��;+$@ӛ���J��V��:���@�)籝x )?���#̒���86b�&��L����~���3�N�d��O�	o��vаS/ґL���֍���[!�� 7.�Q���?! $ω����P*�d8�6��x*�&�l��#,wfe�ͭ@2T�~�*s�r�ar��9���n����šYm���ǀ�������{7�6	C�R��Q�ŸGp�[q@J^�F �`ض��<�$������9\�5��m����u;�z O(\��5�TD^)�n�pփ�f*e5��-��ǃ�
��Є�z�x�S p�,���r��l��S�(v1��8�y���N3a��l�?��g777Þwܦ�ɂ��ْp��� �%瑪�Ęh��SӜ�o葊�ef(�
4UU��<����
�d@`/!&��SoW�����wsL�B�`�3�&L�UBB9���4��Ϊ�A'�>6��7l�Þ��t<H�\O�&�9����NP��feI��-hɂl,A־IP�*a>��I��ո�yC��l�B�w��k5�"���N��T3"���F��,0m��[�L.Us�@r{H�8W怸) �|�}¾�����ח@�Ć�L��gX�iw�w���̊QW.P�@w�^�50�X��l��$Qz!�J�	^g{� VO=\6��Hj�Sj�g�� ?9Ut[��4&����+���%hR��?a��oH��c2w����kU#����|4{SS��Ë�����M�{~��9�r�E]WH�8X޾<*�?����t��Ʒ����D�lll`�5��u4��"E�АC@��Za�qT���m�ܗ��������U�x����$3�A���@OJJ:��GAA!^�]�8�:K�(�5։���0(2TGGG8����v��rS?~�tJ�(��M�q�A�>��	�/]�[B������hC�:��R���4��|%�˰#��Z��s\[�Sؘ}zm@+rb�%,g�kx�����(T�@���밹:��y�啤�JEkw���%����s���M��(p�����uDrF" ����S�wW�RY�,�>���*��	�y`����䤜���o�CQ���LLI�65���1Aŭm���Y������}�uh��MՀe���ct�M0#�, �`���VRu@І���^��￞��c�g�AtT����t==��v�,L��*6��r�uvt,/Ih0���;��G?��Wy�`��d�
F���wVS��F9:�o�c�l����d(K�JK�S{v	^��w.�"�0O��?�}��qkFʜ+a>�@���<����B�tGd��O���5#�࿿E[�?��S�P�@@@@2�;���1c�@XZ�����QV�:{�®��yJ�f�C�f4�1 ���n ���vv�l���с��{-,Y���Iۑ����Tv���.���D�� �R�conJ���ȋ6�O����i�[��b	�l�hnv�GH�#@���723Bwt���C"#����B��antq���ΫW���`y��M�3��}����`A���f��ݻ����qa�o��1&��|2�D�����'��C{:,Ny����$���n7�7\�$r��������
L�ə���8O�Q���l�N�r�><�y��m:[[[y��Ju��o�\J�F��s �	Dr~�- ꖂ>�� E������I)u_
[
�%��	g!!��8nj��/=��<�(ih"`���4ny��W���,W��ç={���"a�������u��x֯��/�}U{�(x�B.I,Htm�o�}S��+�-����[prr&(�WggdQͤe��G��ˉ4-B9�O��s��LZ�	9
rq)��xq���ߚH�
^6����v7-*_K��-*p�z�f%"*�����S��vǉ�HKXo�(���f��>:���R�*)�q&��a�����������7�Ps����{`Y&���qۋ֖�#�H���$xR7�ʯ� jE��)	S��Z�]���:���!d�)���7JS���ɩRڪ��t�#P����p^~v6<81"y�p+�Ed��4���E�(a��l�
b�0�%'?�a�v��k��Le1�N^�j'y��cf��܃;��������JLu����=i�V9��<���]..����]�������z
���M����:]&y�>:�P���&��O�^,((HmAs[w��ո���5d��x��ϗu�����sO2�����)��p	sX��X��cܙ�5��,i�͸�������E�F:��@��`��߶�VQ���������3x�֐7z�rh��.P J������ut�_�>x~L��B���!��].�����R�
=�y���<����]:��j@>u#�G���褤� ș�@���v��4�����j�����]�W�{�܎�NRm
t�Y{k3x�N}��!���^E3�/>}��W����<��C�w�U���Z'��\_�:�`!V�y�(�9��n��۪]߿sE��?��R�R�Ӷ��Ɲf��}D���ҟ�J:9��Ku������X��a��{5[&��H�i��7yv����i�Gw�uv��W��]�!���$�ù���%��QR����ظ'�*�VJ)��(4L��� 
�73�we��a3)U��斖����!@���ě8v�~�TYQR���n�'�7RE�A�		�a��{��H-�+����/c��v� ����+��lfi����aNB���x�Y�]a|��7����hmI�]��9uܞ$�p}?e�q��B� �^bzX�5{�X�ě:�AED�S�9���ER܆~r��̠r�Y�#��x}��pB�}���Y�Z��{yy�sk��l��Ȓ ���Ү�=��Z��xҌ���kj��~��Y� "ஒ8w�|���p�ѣG�+<�0�trU�B�E��Y}]O��a �:i������v]�D�n/o9phV=#   	�}+օ�s������^��Yxq�_�k">���S �ݻaad嘊^�������Z?���WC%�2/fx�b������</�:<ئfAKM�T �-gq�0����n�>�iS��x�b!741����7�E�oL�RWoo����\��/K��Zc��7�?G	țԊ��+S�p\�9�(GB̡���)��׏�@�xFx`�a�x�f�����X����T;��.܏n����2�N�	��Vx3��a�H6U�'N,�XK��xx�wk�'>9-�U�����'���IY�(�A뙖S�0ޕ��)��툩���Q�?o��Lś~��s��bu_�8$z5�0e��v{�oa���"/>h�9��7fe-�n�0U�%�<�?�l:VLL�k������\�n�������m�Ǐ������*w*�����t��~���ƼZ�
H�'oq��~�b�6�dr�U�s55صr}^��B��
�� �m���;�����?y�<#6������}==��"�f_"K�� 9"�� �]����;�o�,ː��� `�C���>�����?�P���Y8���D�)�ՄE��*����ߟ��P((,�����N�F���.�/�;�����=���� +n�:{WJI)\�]<l(��;
��$��:�'ta��Lq��� �.V�P�3�M�vu�g��q��.`����H�j�e�"CE�=�(�d��Z�}tIᅾϏ�$��c'�@qXM����<��.\]_�z�����~xGo����__pg0�ncw�D	0B	2�e�j�[5�7�.
>������@�I7`�8chkKKˤ�� )p�[Bx���͙�����mnn}'J�W�6��S �`T�϶� N ���
����{�+m��ۺ�x�z�(����W��]�^:Uz7�-�e`$M1�L��b`PZ���\b*���4g��� ir����;u�>%��Ǚ�ޙ�R�vV����TD+\'�p��+^D���bk��)p�\��������_��)�ED2��!���A���%�Η�ݼw/��Tz^7�G!�	�m\Q�F��O�p!U%e�����������N4�N�����#�nth8���K���ږ�-P�o�8��,��i���p�Z%GL���3P�upU�\@\��-�V�S}�^���׵�"��\	�5���1lX�{m� �ce�!LA .�2G�5]T��V�?�8O�C	Pr��[��*y�x�{)�%ʉ��TD-�}�7�o��RS�Ţ���?�n���}�SKu��x�jhh��~�Ju1�+1EJ�?��&��pW�5�d&�]��;�FYP@ ��ة��ʪ2(���XZ���Lii�@y���-:"��}H�b��
���C�k��=�]>�u��U�2/�P�r��I�S������\��Dg���M��n���<�&���X�Y��J;k��{��*�������$
�,�����9���ةd�|8��=S�ڠ4JRT�Pmo�W��YPp<��M�VS�Px�� �W�_f+99;-mD��0	���'.�_�(3#;�-��Փ����}n�I؆������e���֖&Hh;��"y.aᑙy�L'�U��u�Ā�%���r�|���{Y.�\&����kz �3��H[����E�s�T �
2��p�E����1h� Z�]�=�k���c�:]kZ˷#�ayd����I�uܮHׅ'��	0iBZ�+�s/@������d���&��Mx��U-��f��G�]�mw46���qT�gan.��)b�G��=�^5���H�k��>�`222z9ڎ��>\�[j�c�~�Kl�}7c8k�>����N,g��t~Jd3���t���qd
HZ�|�.ћP#�K�%�yDx-'ޢ��-y��y8����q�)k@!���@AU��X�0~�?�llmq�p��[Yɛ8o�їj������t�Y �?�n�/�Ǚtؒ�����:���%!qₙ�3���ըѓ��
�����y�iDN-���3`"�]��}PO���+A<�״������&9o��\~r- 	e�% J�eIKXhd���ؙa��չw/�D�zz{�3'΅��g'O�4N�`��36K�I����H���_��n��i�9.� g�uf@�z�$x_�WB��lwҡ�((�p��Ny�=����P( ��9��l|=��V��o��|kzA��^@��$e~�����J�vNN���f��"����y��7�{S�͐v(���������X�ۗ�2�>��{G��`j� !�}+�=�U/r�`q�؟aƑv;�����R�|ݗ�O232��m��/�N_�=�����ܠ�r���.�=uxE?\�'m��d��t~��I��c!l�	KA�T0Y��cߎi������8g��yA���L窢��Ʈ"5�[JCtj�k�`C��+�X��.-���Z)�NJ��:��i�Ǽm�H~��dR�7�y�s6�c9�:W���l��)��X̼$���6�ޮo�p�v�@)MF��EN��M�L4Qhe;Qi?��q^Z����:��p���t���LO"���:T����/w���hB��8ߨ��w��#\d>`|Ht?�t�H#x^>7����;N�����)<��uoE�e�m��M�=�����4ob����� .�ܖ)6�L.�q��wa�)XO�Og�*ކr�R;�8� �x���
o�Y�3�Ӧ�����݉d�8��k��LRF�e��`�%h�5�q�mi���%�fx�-��w�fy�Ny�@����.��>zJ�m��C��������c��u:]��y��+(������_3���y�Z���V�
�@o�S�.7i�w�>L�b�;K�©�.S''M��|%���}ܗ�*��*KX�����n&�^Kg� �f��Y�`o[�������А|�Q)2%��$��QS����ei�'P�����!�7;�,#�[�DS���n��Z-]b�ac��(%���%�аo.91^����x}�Bn���Y�q� �;
i/)��UP\\�.�H��3�KZ��uOa�4��L��������H};���v�y��Wr�ovx��\�u^����@|9�����W�c�kN���~��&����R_�:��-U{�b?"��V{u�|1��L1�}���9,OPl�ޜ�S
��<~�{a-�&����
��@���+����,u�e��<*�ϟ��`E23�f�}I�������,�7g��f���+�q����JI�a�������1���y`��[�Oxδպ�o�Ej�L=Un94�����:%�׬<��ʂ���pB���u�pXꩮ���IĤi�0����,hr 5�ùp�M���->���5>;K>ߘ��GX���zkA��-q�� D�پ�F`��C����|L��C��ڲ����?ќ��E�������|�~�2���L�o�}�x�ʊ.T�|��="[bWI��.��2��h²`h���4�)Nbd�����9��k;���
uģ�+����ƅ�m@���h���h�2�S�K�^~�K��('#���1h�J8�:j;Ѻ�ϙ"g8k�x]~db��}���nj�F��{�(9󍏢�$T����G������hh���3^�:��q��8�YnE�s��;�:%Ә_�jH7���\���Y��}��W�ښ�A���+�N�Rv[��G�G]��-�ҵL&�ŉގ����ץ�f����@���6c��DV��6�p')g��$���O,�B@M�E�E�����,���{�إ���5���Dl*G.�^��N+\��_s���
�y��W��NnPj
��UW���7��O#fbzJA��z{{S�"�vZ���Ɋ�	ҽ<�a 6����]p};%P}/P��f��hM��.�����������;�Zw�������H���PGzwlt����%)JJJ��� ^�@?0���H#�V�=I���y��d��S���YUKJ�L�1�vH��n۵�򰮺�D�9l��c^��yė�����*5�.=��j矤�X��L�1A��x���=�2���%�=����=��}鸹�~\�;��cw���|جi�K�f	��+���%�����)9>XXX��U��j�މ����g�U����5������U���GyTDi~q��jͼ�[7��5���hPѭ�w���"�{v��az��b�9��� B<��v)�cB�^��>?��o-45vr�YMY����)Z;zj�}"�KW�j�&��p^ρy�D��
Fo�X.Bq���0��-,,�wV��mx�<v>ƎN�w�Ϲ
�ib~���.�|撮�>82��!w��s�i��ް��w�Uh�H�knV6��pdd_�OήMu�E�İ�Q�������lNV1��n��������g����G�t) ��[��8��_Pz#`� �PeL�`�����y]�rF�I��q^��=���#f,��
)@hwaY8|iq�ÖS:��wm�P2�2}s�� :�ݴ#�t�!��;𳟷�q7�Ð�v�8�-r];J�!�X�V����1ج���LڈYd�����6��<2���5�#J%X{�h��D��E��e{T��ǳ_?	�07b�8#M�
d���Zx$�t����̾πzش����gn�9wLʷ[� TϜ@���Ё�p�w�k��F��w���a*rd�%%�"�P�7�5 r��Uk�,(� ��ί�dK8����r�V�sGE��&1�LʙECb9g��jR8�_^^���Ao�ϴ=�|?K�9Z�h�S�1���W���-+S�:|�h���{c"�f���䮴΀Ä�n��vb���u|8'5�G+w���	T�;{�5�:���t4�k�\7yID�02�*t1+�=�wN(���Z�9�
j
:��>J�#޳����xy�ʤa}��vI��q*X^���&�^\& z���?U1�q�p%��� ��;R���[���M���KSS�Sѽ�SB���R�L��D�n���!WF�ܢS `��M��&5�+���!��Pk	���d�����'�|s��d�������h�Z�����
�v~�����M�%TO������ƥ|·k9������"V��Y������k���&l6mm��گ� ��k�l3��"ĥ�3ei/m����W6��;,;����d=��srD*Gr��>2.t���m���6ʄYa4�(��^΍3 �NC��C6u'���=
���Ԁ]D�����O�4JVT\Q-��FNE��$�%��'�vF7�[���򝮻���5��l%F�h�����mșX��PLFp6m+���l~4���X��A9����n\T\�H����؎�\^$��+�� �AK�Ӯ�1=�ZwML�&�8[���2��Q8J�Do����*��!��'��vE�bI�<��c��*����X	P��q~I8>N�'�~qP3��ʌ%�]������?��m�ck�U�����GAxM�SAfdui���W'@�aU3==U��R�_�����+��jY,�@b�GN,�?���>��K�9h x�ǫJr4������ ˷���ù'_5#�Ăv�:�H�T�8��F4�Eڅ�cҥ�Uޭ��ui�iU^�/ɤ9��i�H�4ƕ��mh�Ի��3����N"�?)L��]��N�YwjB�}Me��)�mMV�Kh�É�BtTQ�q�4��.>�Ǥ���jy�y�a��Q��~�|�Փ��>�beN�Ҋ�!��>ڼ.����N�wp���	t��O�m5s�o�}:N�$$$��ke:5��I�P[���l��OT,)�+�쵣�+�;���~��!�;c����*NX��H�6T��o�V;�R���0-\��7��Kk�;4N��{�,�W�x�v��q�*}(�.0)&*���^V}f��\53�ro��� �l%Z��"�y����*�Özz���cDE�:)}�LyN������bޛ<����Y��uQ[c�?�;��n9�#k;y��ऺ��PSt]+�l����Gw��	��"ҟ�(��&a��ҧ���|��FjZZ�f�X�r��7�9���WŉQg�ͦ�T3yA])��C7!���s�?��$p6�7�$\��dZc�Y��f�7FI쩣r����Ms�[8r�|X,�-�;����Yj�˦xR&Vy6s;Ǖf��p�{��G;�"_ol��_Z����﬷�$����2�7� R� �xr���%=�X�z�Nգ�B�E�]�0>~׿�=��]�E$��Ǯ�q	�;��}:&��V�[	�}:a⇎(�S���N�c��?働w��TQ1�^����wz�,_����uj �#�4�T:9Z�;���:�7�#x��}����V���=w<5���_r��{7���j���:�ެ?X����ꎷ,~?�{Hg0�:vv���%ed�����S+
�6�N�&�in�i`�V���f��{.Nff/�R�Lу˾>��ۦ	�;�jc�M�+�k��?��ʖ�]P����]�:���B�irθ�.j-��rV�j|��S An��Z�~�TB�kN�B��ǰB6�N-l�T�͓@����4��+B����l �'���{�>0* x2:�����4�Tj�̛��^[���`K��@pP�pٲr�f��p��1:B�:A�kdc2��k55@,�[#�-�{w����׻�[v��Hr͏�q��x�c�7�ۂʤqKns�L=��:>�\��e����\]�ol�@�y��̄������F�&ϩ*X�����/0)��@II�h�(�<6� ���Th�_� �1�Q7�W �r��{�<��q@x�ci���$��ᵙ��KB�4Z��16�߮�����Aϙ27JT�q��1INΗ����*��4)wYDb�^5�w,X�ϧ�
 ����a�Qt�Ph���/�7�Sy��
�6�uX��P��n+��k%���y��@ ��}�J)G�x�UT D=N��v�Z�K�L�{մ�۹Ԙ&�7�)�bU�=���֙�~���s�R3�FJBJ�ry߳Q6�+�/��6�s<ѓ��;�M�K�(��>h
u��,"z��<zP�w)Hnqq]TPP��<��wc�\��[� ���V��������{�I?.��JĽ��SW�bn�*}>��2�ju�c�:�ز��L�&�Ǽ~O��ỴTiP3��s��d"$՚2j�ey�{��D�Ǔ��~9�M8��)Hߝ���y9�	���ڭ��� ��|���i���c�a��"6e�6A��3A��)����e�]�+���~��/���㌝4NZ��q�㽮$ ǁ���b�vݸ�<&&F)�	I��7���`z0Ѳ�LB11~���>�6y���͠���B�Dtx+����We����V@vL��L�r��).�:���$(`#,4�j�۟��Ȳ	��s�M�n�=����@_��:0�9�G��'VդiI�Y�(�y ������b�5�$g �h�L�}�"V���<ш�'ml�q�S�];'�A`���R���~�+s[��+[a^��%P�ɤ86�t<���SZ��U"r��m�*�T�2�1����#4�:w����M�;��M`JUS�".	�׃�3gSTN\'�YMv0��
t�0��8����SX��55��F��0w��I�>�$A|��B�
�h�kvȠ�e+ErS�|VL���7gu���xc	�R�Mic�R�ȝz:���E�
�T�n������`��uB���f�Fᝡ�	�aa}!�G��y)���NRr/k������D������_�;����WO"��)WO���ea;jw;��8]�-��t�V�tdܯ�<�-�s5��T`Wە~ms�|8�\��ƅ�#�+�5U�r������IqM�Ud»���-��5N����!0�iHI�1f�Z��7���t����^���^�O�v�N4mV��T;��6W5��(B����'f�#ɏg�;f�i�@U[@�%Xp�Z���(XˡI���Q��嚨W?3ip���H4Qv0)B;J^�c␉hRw�S��|ٚ����b~�n�`�v D=;1c��c��<�Z[��vWr�'��?>jx�����gР�Nn�m�� �iH�hP>�����B��2?�Pnd���f9x=�.�9L
X�ϟ� ���7�ZW�m�ԍ�fi��nK8�b[&?{���/�W2��Ϊ21��c�:��0����2?�ML�
םu�S\t�e<��᳥������"��~�j9Nd��e�>��.,�AA�<�]�rp�<�PD��������r�{@ȁ�G�(��-����|�����}���K��yi�/�, n3�B��_�Z�<�m�y��05������.k�Y_��6��.6�h�]b�������Lf_�;p۱r�bĬOg�2�R��:��re�1������, :D�L3�T�o$���IX"ߨ�Y}E�3WE� Q'�m����l����$	} �p��-겞wYC�����.3�?3����擙��(
�OW8��J���ރ3Q� �r��,��,�/W�.Z�w2��_x9s|��l/e���5�RB֧O�s5�U.Yq���G)��m��:�p=թryVQ?T<X����S(�s�G�E�y4p��C\���"gl�/��=�?֎W <�hQ9fe=��eh����1��0��n�$�O�B 4y���G�^�=)O&��J�І�������v��u<�2A<��Х��k�h��?�M�Ϟ���??�Wcǅj�=nI�x�����qԯ��I�5�.�2�a}&?� N%�S����)2ip������EM�g>���K�a}��a4�E�1��z�?��k��߫��+캨�|�.�䯨��SgD]�E\c��q�R�qi������ꣾ�*<Y�U���t�|n9��c�oK3�.k���VW�~��9�H�-�����k�z��W}�1���]f�.mB�8����Wz\e<1���_�1�7��R\A���X���>�	�%X9��Kf�69�3�_s
������I�V��%�G��U�s��l��c�<	��Շ���T�g�I)̾�#$�m��2�sg`Щ��Bׇ�xΧQ�L�?���,�#Ż!�W�r�y��LB->bQ�����cʋUk��68�'{�#�c{&`���S�3�x�����t����Me��)�@��C,>�����KXy��ņ�pdx���³��N�ɕE]:^�j���Q�[ W�Xz�69��T��ׯ��N�~��/�.jd�U�:�(�]B t2���i>�9|�:�g�c �ߩ_yԏ�dSm�GE����X��&�y�
��X 8_�H�O���!<F,�� z����r�k�qTG�w_^'�jh���<A:��j)ـ{]�FE���p�u�[���S�Y�ƣ2kE]]D>�m�@�-�[g�?ġ���#���1gT�6E�/���Y��|�����vr�̈��A(��+�幊〕��%��@�¤i`?V�s��`��Oڛw��(���D���W�T�Y�@{A u��ʄ�1\�=�l�YqlB.�O<�h��@_{�C\q�(p������~;]���������>�whO�q�sY"o��/V�A�Q�#����L'�>���g�
!|�Ņ�h�1������ �d8u#�߄�~�mHqq�}�P�go���������K��]��q�{�8���$���{���i�Z z�3�=�v���*|ĥl�r:�#VBj���q�Q�x08��Yٹ�!�H�qY�l����H<��4f�', x�=Nڗq�YL:��ε4Pc4��8�z�W'��?P�k{��#�F,��PGm&HX�zL�ћu-�[�擘�{yEY8��8�"G���������u|�0M <:s�"���,�2�׿N�������c5�Ï��q�0Lu�[T�(/`la����S�h �KT�9;���*d"И��V^��w8���o���i�T��c�n��:;��]�#
���m+������bb>�)k��_U_����J���B� !k�,�Ⱦ�Ⱦg��8E��ًP��5[YFckc�a�u����:�>��9�3�>����u_�u?����˨?2�p<���@�j�`)�*ႚK��)ϼ=�'x�AWu���xO��;91d���e�?	�R�9#��Z���B�w�PA'��E���0u��bD�N�����yg��hP�4��L��w��"��2H:i���0�e��z�{A��h��66�-�nn�%��s�9��tN��yG�PA���/g�P��u#d\���d4��x>'d�!�W��6�Ss��G��~x��IG�~�ls��Z)߼bX���vJ0����с9�/6���0�S�[X�P�J�]��1�6��[��u���������3��Y�wJ~X�3I#�����Φ�2+�����o�ܧV�;��`�O"�S��$���s\���RO̓\N�i0H�΅z�@��_!4�Ծ��.��3�ڊ2�T�T �|��|�EMp�� ���)��7~�{��;����� 7�������W*v�4cq7����;��drԧ�����������������$0:�a4B�3=�[,.����/���E��z�PKܩg��u����>�}�Dx^Sзi�����[�2#u����@V�:�89.�'��/h]	��!���N5���k

m�E�� ��<ʹ�"�Jp����T���ɬ�|�sYa��>��bW}��=9�v�ʩ��%#>=cqpMD
E7P6��]�w᫥*έ��h<�Wd=b�c�ؚ��z��~@���+�t�)��g��A�W��%.24fG���5���Նw����ӍX�$�PP�`��՛.��R?���^vF�8��� i�7u-�,WNVYV���:�s�2��56�'�����|�<S�|S�5N�~�-���������I���*�9E�c�sƄ�z���U ��U;�b�J9�n��Wl	%����8��x^pg���6�՛�c�z��n�4��ĥ}�h�QA�����Y�e=�, �b~����y���g��25)h���W����T`)�������}La��,�u��zޱ4��K�fdN"����N9/��a�3X�K%(���0��r�;��X��XY�����'��t%gf<�"a�gV�������P�6X��+h�� g#W�_�#T{����Z�@�l����zKS!�h������b5���kD������2O*���xz	�:��p��_7���û�[~�g��-�e:�Xb,� Z�8�nq�	��1*OuDK��O8�loE,7B�C'\ezS:�rm��Gy��1�y3͔��I<e������^������Fd��rm��v��!6���Sc���<��/{j~q���F��/LʼKwpE�+��}7*�%�nt]"|{��?d��)`��9�J.d�0�o�;>��3���@~��'\)�(�>������8B<F).Ru��v�ֹ/���'��	+;��QӔ:{bVW�W�j��6��J���tA@�{w�.1��:�q!�w�X�m���o̩(��2�,W
i�9���$�Mo�:e.F�;8��Ӎ���E�?I���L(n\δ�x�Y����W�����Qi���� FӖt2�ʟ���Z�(�սV��x?K^]��oL�l���wa>���d��w�x��Αڑt�5y���O��s�T�e/��d뵈e��.b�N?�	s�G0�]V�љ�q��"+����@�κ,�&Ԍ�[���� �|�4�D����G��Sl��)���:o6����v%j��c�a� ��P�^Y!�H��&z.N�'�и����27Q�j~S�u�L�G_�.�D1��I+p���w�9���u4/�?7�i���b��"�	�Wa;��<����r�����j˷���y%ɧ���W��sB��~0��~��A��O x�����,9�{S�ohHO����⢤��9����2.r[����{^�ݜ��m�qC��/E�:F�OG��ΘE��4P������_R�-��QY*������o�r��fM�]R�q�3�o�_C@THX8��^$-s�.с�s؇C������{)���5Y0	�N�k��J�E�z�DOdD���`�a ��-�7<ML���*�ϊ�h���h�ϔi�����>�[>��ܜ5fbK��U|o�ݖ�5�m���p�Kk��Z|E8��+��6�ֻRř_���>>;�S����d>	�v1���b<D8i�D��muT������k���~N?I�ʢ<����d�6�_����ه�wR"᷾���5dY�ץ����0��\*���ZC� �-Lڪs�uT��N��i�b�qk\s��r�-�&|� ��؊_ed�ѫ���W�����W��_X6@0�����J>�5��B��� N�o�E��/�hI[��x�a�I�mj�pG6�;�5�͎���	�9���@��Z���b�~K��cLT�Z�#G۴�T��lQL|��U3.��M�ٝ�;sqĩ`��'��!�s
�gG�'�I���3�6X"nٗ�:k�n6�5�rR�È��RN���G���K|z����1S&k$��~^>�>������,W��<�h"!��tQh+(i45:uq
T�셨�(m����~���:2_7�[ȩ���Z�I�`Y|��}e�����10i��,�t�/�����rP:�j�f�g����}�[ҿ�zPP4qt;�)#��SY�Op��������-;'� �l׫w�x�Nڊe�8nԻ�l���]��[���6�����D��ّ��蝥���Kػ��9�%��o5 ��t���T�d�1%�
���qJ�S;W?eU�$����E[)��+W�&���:-�e7����3���l���ضsh�{�tP��J6WE�4d<�\�|�/\��DuU����	W�5e#�y	����f����Z����!*��lU����G}��M?�mL��}y����UF�T�'���#n� *6(� ��".,2S�Vk���ʪ�x�v��2"�n�+.�'�NSA+�V.OƝ���1�Kj/�/+��ײ[�c���w�p��k�\�FG4y8��is ��YVᮠ o/��3ZJ9�xMw ��!�{.��i!����c~�w���-�7�}�v7m���ܞzxm�T޻3�M�r�'C����G�����a���B���m����K��4I|�������c������8Ş>9��k�y(��۬W����~Q+qת7�P�����|�+R͓~ȈT�`�IS��DBm�Z�5�UpE��7��Tl!�	ヤ��n�o�P���C#�_�u��h���G�(?zם�a��J�7�֪	S��T����3�� �p�-]�g�{�OF��>y�4���{�����z
jp��fO����2��S���<%'/����$5*�/��]*l�N{���+^��� n|��!f>x"Gt�]�V���;�Qߔ7u5�, n�	^[�S!B�7弓�KBV������weE��0t��4l�Uo�,#'ѷ@�����̷T�Oޔg��]���'*$����taf.!� ��o�@�k%>���F=��B&m%I�)�z�ŉf���=8؅�n��K4n��IR!���T�I��l��]mp�>@߸�B����Sb�J1̛���W]SzgTT5����,Ƣ�MH�7�J-�/SrrgΜ�a8Xc(��}XT\��s]ހ	���6����ѿ5��@K�x5�-��{s�HvSTM�x�Q�p���U,�4B��|�;�����E>笰�*�k�:ou��$(���jsޤ���wr6�X�ߑ�I��ז���۾z;����G�2@I2(�qz�y�E�m����Ȉ�x����Q����m�`?J���z�?��K��-���;��$���%��¸v���De�3!��6r@A�7�<��/K���|r_�R^�z��MQQ&�e�7]P���N���]Kw��%͙ż�(���%�'7_�\�2�OW Y���p��s�gם����J�,��>�3�qrM����-h$ZňQAkW~� 1�7��ϒ6���>G�;1������,늷v�4�? `��*�w|;����n8���.���w�灄�������M/P<.�oԸ��C�y�U��&�z�8�����<M�aNW �-Ҵ�d��ٗ5hOG�?���F�Z� 8��dE�k��%���?�6"Hr�s x���:��B�$��|��=���Tx
�FuٚH���)5�l����5�`:D~�tV:`�{�E��Ē�����	�\ml˸�O�%	�ܚ@��o5L��Ֆ8m̬�_������nc&GT�$��"��}���׷����|��S雪"aDhs�Ff�rw��s@��L��`�Rt^a`Ǜ����Ԯ�W�N} Y�_3�����*���t=��¸y�{�K�����J��4��LMo���:>`_9#8+1�= !����Y��I+�D��i���݂����_t<����}������g	z�K4M|)ڃ+E�2��`�lԛk�=����f�0���Ulk���!6?��W�+���I�C\�S�,?��<����*`mcC����T��`���>��љ����L�հpM�Ŷã<��KE2�md� �~+�lV��g@nҗ�Y������ʫc�#'������Q{A_���@�H��FJ�8� ���,�.�[n�"1M���-ʴ�UQ��\��\�g��ܣe�KK����N��&Z��}�َ�߉�9����]vk�)R�ҸS�ʕ��	��D���m���(���A��s=���3���v�$��ʋ���Mou��+n3*0�|�ș�ە��-A�>����g4d=����� {e�~A���4�D@�����w���?�7�!O��߯��p�M�̶r��-�nS�O%]�n��m003����t��RKLL���pVmN#��sI]�j�z�/�J$�u5�i��~G��h�a_Q7	*1s���pe�z�w��W��f|�� NI�=,�����n 6���&�
XTv�2���w����%���+�KTé�?�u�O12n�
g�be��ʄ�Ɇ��)T���T��5�a��Hp���J�f6�ݥ��V�K~^~�+��ܬ��2��t���?��{ȭ�`��j��I*�����/C�&Am����ƺ��C@��{�6�u�$�"BqQ`�^A����NF^cMj�ďg%�39q�����V+�Ͷ���-K�V׎�}A�#�gZ�gR*��f��>Z�J?BЙa2��W�Ć��Yu��!���J��6U*޷o跈���V����S(>�]����$ ���$�^��ד2p'O������J$��q̲FǢV;����V����C;3��=S�� �aQ����߃z7���X�� ��_�8������k���yq��\ҁ�)���q��(��!�Y�-�+���f�a�Ԗ���̲d�D�U��_`r�P���0#�\�x-*��؍\]�^���d�����\��k��f�t��'㺥>��Z��L���awc�.�9��l�W]~^;Hfw�NuK�7�5`�Ь�2˩ME�)���x'���r÷vu�:P��S����b56��	q�t���e$<�L�E+���C�b��v����(�O��?��L(<�ߔ��+ �7mŜwi�Xٙ�Yj���"�Zu)���wi�����O�y�D#��yD\�_d�z�R��gOµtuK���N�p$��?LTir��K���g��S������6T~�f�l��H�B��NG�&�r�����P���%H����}a� �k���Zf�G*9:9��b���b�����l�=:���SQ>o������a��e@��"*ME��2+���Y[/oܩ�%;z.oX��IWU��<Ywu;6|`J���"x
�*"�������4Y�Ms��H�_)_����~v�m�6 ���W�ў
�'�z�Fj�)��*"��׈c��R>����-�B)XM7w������.*��Ld%��c�ڣ�������RZi�2o���ժ��Izǰr"�� ^�`�ٶê��Tu݁��;1�����h/ח��TsY�u�n�V��t$<��wwhl�L߄��p>j��^�]f$>���t`�h�Bƀ�J�Ď!{d\.��
��3�͑��$�ک�8���Tj�B�)ߟ��%�MG���s��i�iV�c���I?�Er��ǳ��O˳݈3�[Jm�K���Vv"�eu�}�ƌ�_Ʈ�ɲzY\U��l��ĝ0�wĉl�L,&��m��[$�%�����f�O�2��D�����_�"˄$��6�o�ڊ�/m��_�)U�i����,�r��d�
�����TA����r��b�ڽe�d��MK\L>�e�@�na�۸'�]�*
<�2��U6#OzSOck�ܽ��3XRҕv	,(E�����g���e���voS�S�9�I.�:���s�-���>3�T����{u��Cy9
�r#��F�ӊ�q�V�<�՝�����x��فE��q*=֢�V P��AdE(e�×�����+�n\u��X���<�e�jGJM�j�Ow��|M�0#G�0�/��א���ɍ(���P�P����A�{&�L2��l��8��B�nJl1w-B	@͹]eB�v`����~�֯�74LtR�y��{�<}������P�qhʺ��~�;`fMf����xk@K+x��Z�Hߺm�D�`�e�q��C��G�����d\A��J��y�gD&6�.��$���
e��~�A���,0���ībf��l$���+P,)���ѽ.s.�cԅ�oZb����V���T:,��JbX �� �Ě88r���5L���;�����`���Ck���*�v4䘰�./��%f�Eg�&���}fQd��%I��ɆG�����^��&�_1�9|�`ȟ�����Rh�8^�@Uq;����Ŵ�O�R� Y  � ���������سp,1�(��%�іR�z�h�o���ɉȵ�b�k�g؎�E�b���9���;W�no�IC�����>g` %�"G�u©_<�s�)1^�2/�( �~[fee�~�K554޶�5K��玟i�e$�P���
��W����>8��r���������)l��T(���m�ba`-0�A��E#�(M�E�M)�O�1�!�jU����]4�;��\0��U���u���������8��Y�	�`8�(�KW��AfS�~�53]]���
�BCn�q�M��W-�<�ޝ2��bKS�l��z�$���[6�������N
~�M�� iER�*b � V.��JU�D6q�\��ܜ�DF�%ZU	�㛕����$�we�D�(��tZ� W�����b��W�֮�6d�xAAGR���g ��=������Z���=��yU��A<�����n��~2tB+�
����܌mX5�ܒ�N��:AӰ=ŗ�ܑhl i|9;�O p�}�ng`f@e#S� �#*�
�����"���F�L-́C8��`ZItO-�i8�!9�ZsFq����a~���Cgʯ�ѽ>D;nh�齗��������� fY��;���byA�c���C|.�m0=y4X��&��[�<����k��N���h�qI�H��ϼ�[����@�
�#B� ;�A�`Z�m|�LL5�ݬ��Xꗳ����rg?��� P3� P3�:���j��瑝�Ó�Q�>}��D^���x��C�އ5Nh�8h%p�5����ݎ��>�|�7�r v�����Bd����P*�T0��8)�p@��=('��q�Q�X䈣%����xU<P��&������l�-��X�Ȥ���ל��'oPdNsz�մ��}�݁�ؿ�8�]���2!X5MO�I�� �#{�^�`0l���̊���җK0����&I��%�#D�U��[*�;�G�kvv������H<�b��o���N�X���S�Hߛr���(�"#�=L���I*}2������Z��_�e�4��G,��f9���['?�FўB�T%&�bD�Ŋr_��}��M�&�0Q޵��U�{Ǡҿ�s�EEG� /zH�wÝ��F�#=��]ř����oSCS��8������͙�]m�2ҁ���)��F�������<�ӥ ��!n̭�_nCAt�v@��V%p�FuβE*%��S�O�� Ã��U�ʥ� N�>o����.�����e{(g�T�|4;4�?�ݮ�L���yD��~���1F��xUf��x��չ�h7V�y6���'H�����t������]����ce8;��cRD���ll�G�b��]K>P�f��^��X���r���H�?�����J3�����Y�� ����ZO@�b;�\E�i��3��S�_>B(��1��&w���))�w	 ��ln'��ۥt|�����l�[�	��>%�tH�����_��<��O����Z[[�N�3�a��� �0����t/��o6z0���~�~��(�8i�	�	'����S&���%ݍ�,��v^���Ŵ�J
/��P� ��>��I�Y��=S�Z�Y�	���݁��]���F.1�B
{Q��?���AJ�V�p��D)�04JIH�?���t���s�
*m�Δ��A�ӛ�i_�M�nNM���GH��Y2&r0`Y*��Q�2�}rW4�Dnt�v��]�3������=�œ)�]���� k�K��� N
e��̰Om�������r�žr�)�e�?�}�h_�qv�U[����vtQM-Vz��0��`�R��>+�n_	�%l����<A�擡��0����X��=��Ȳ2��9�I�z���/� �p7� �0U�� 6)yz��(H%�����om�^.YY�T�j�򣤜\ԈcU�j_���nG3V���D�ěQB��6��׃0�&����ڞ�*��"5��.u����A(6���f���%�)��[�kr�P��1(�<O��!W�z*�D����yz�����������f�j��ɕ�u�`z�6$]/���;ܒ�����p��fQ<˵��U�����^�gb���zX&�7/�@K�����Ez�eB�] D���LMw�J�0�j�5
c3���VɍC��cx`�Ez((�� ��>S�d�Ҏ�q�f��"�;�j�� ��½ `��]Qq�*�V�_2�l*���@�%�k����}8���/��Vȟ�(���m��.�T4-���\��x�8^��v�@��l=�D��+��SS/9$pZ����ӌ��!����1 ���B���_4�0��sĲ��� �=��@z��T&A㟀<�+��X�
�h����|���+3��u�x�fCT��ޓR��c��

����訑j�ƈ�:=�w�} >ک�20��s��cRT� �,��W��lB�x�fk�R�zׅː�G2ϟ�p��� ���>Z #q}�f����_i�
lĔ^�O��?~��@Fד�|a �8 )>��PG'�����?]s�j�ss
 'C�@�ۊm�٥(�&�>���:� �RrO�!�S�i s+�ڴ�㏞~o�w+PCA���2��u�m��10�x� �^�����k͹.����M�.�����(�H4������8N/Ӈ��x��;�5�@0��O/[���%HI�̊��U�J}*{�M��I�C��&�I��l�j�tu����>� ��&&Kv�9B(����u�����z��g_WM8���[}���'O��<q~�a�tT �aW�9���kZS�sߧ���&Z�����\Gy��=mfE� rVd��wcO/��ˀD>��h��.�H�d�xs]�z޽��b\�yK�b
U�>k�& D�mŚ'd>R7Q,�Ь���o�I�@�eB���xL`SS<]	�e�pmo�
9@Gk��e&]o��$�(|�(,������]Q�U:­D+��
��]#
���Hn@�
��Ձ�����&4���5}��-x���R���+�z���|�����a=�z��Oq@�:�x@2��JzZm`ڗ �j��0/�]�5վҨ	�` ��to�C����6�i�WXɕ�H���䂂"_Z�ͷl��zJ
����i�������K�Vм\�0��)�=�8�P�uA��+;���)j�s����|`x�\���e�c�3�R^b+�����#yf^/�*U���{\�~|�-�e��ԅ�/�q�a3ݺ6SK�n9�)�1%X�φ;\/R�� ���,�no�����u�b�b�_�D�nH�'@�[;#X,�2�S\�4d�
������$�(xs?V\ި�'�����qy�*\;���P���>3�ɧvu��n�r�
M(�?+=%TJ�wٽ�D50�X�ZB�o�)Z�\d`��
}�*H���ד� ��bAA���b�(� �qP�/;?�Z�Ne(옜4M�F\Y��y�JZ�@"�&����0�m+r�XS�3@_�.V�ԁS��[���''3"E����p14g�# �  ����V뎃���`���x�c��'���2{&��k�mL&|�e �� 59��K#�p�S��X�ڡO]� �e@l�<�ܷ!�)vH����Z@�� ?n8)*�Dٗh����/J��X>�ZmD-I���+0��> ��/�I�[�[��� ����U��O˔v����X�B��&Q)�(
�	�8<2�^��{�\C���,�#�#oN�)�K�� �zc��M�Etӎ@���\���Am��ZGq�5�������D\�~��C�c�Õ����9����q��9+�}����ӆ]b����B�!|��n��?��M�en������	�w���ǜ�u���tS����m�r�+A0� �R�`r�k~u�!�=�<3Y����58Ο�s7#[B��TԬ��>��+��B��5�8���8�:]
?aI♑e���Pޢa��4$)�@�X�����N��5���ܸPs�{�����`���	���2��wEz�y2�|����`2k}��*�<g�rJ�?����ӽ]\V�*���K�kٽ\3��΅������W>9 d��"�k�.��,1����<�k��Ԇ����mP�O2�;cOV���K�����=Y7'���^��=���,?���d�%�055��ſ��0G��{:"ѡ\��<o�t~L牖�a���
E�s/ך��>�V/]2���_ݢ������,3�W������ �}{mhhh�a��N2���Ճ-dߤ+wQ ����'z���Z���.ۓ �:��c�<]�&]%�����%����\����r5O�@eOn������x>���'`��b���ַ���#Bw����]X�W@V-��;��N2{'u2����;���/� ����8F�b1ݟk���]�?/��D��<�Ա�O���o ��/2*ڤ�2tQoz���*h�("T#�j�8�G�q�"o閎������cq���q���y����P��D�69t[�0�)䂍|��Գ��78�����n�ED�����^��yF?+Ì�Љ�WȣR�d${׾l�b4-Qh+g$� ��ʮ�0<�k19�WEQ]����?�PK   �I�X
V+c  �     jsons/user_defined.json��]O�8���h���8��+6wlYu�hA@ٕV�r��i&S!��:3(8c�w$q������0m�v�?]-m�5�EY�|:�~�Ͳ�+� '8wg�ʺ����?ۋ���{���SJ&5u}���뺹w�GUk�ʶ���\ܔ��rz5[{z��Bϗv6-ݟS�
JM!�<C�Z����s04ӹ�?O��.MS.��<��]s��\p@�)0bZI�Ɍ!U���I�Hյ{oQVGUQO������\.���C=w�:%�0%ܠ�'g�]�`��fEVU�m嬫���mܗvK���e7�O�SS*X�˃��ԍ{k��6+�s�����;zI�>���!�����o���ݙ]�v�:	��`u6y���脊��4��幗W��Y /�/�v��@>,�zy�[^�r����d�|ȫ����G�R������� ��7�'��B���;��^N/ЍDBB�a8���HA�0�������!�0�_� C,w��p��3I@2�!O1��C�1�<� ��d2�d~�[8$�	/�?:$D������%��!!�l��OB��?GlB��_%a����H��b1�f[����6!�����DlB�寊��h5�|݁H� =H�1�x��x��g�A|��g�S���M��/R@iO�:�Cl��S�ǐN<�*M{��ʉ�<B�)�c'���N����1t��~&T��b�A��]Y�S�� N<Ɒ	'c'��.j��Gϋ����l�I���j�m�r}JwCJSW��0��HVp�Y�#�ARs�.%�:�J�Oæ�]ԕ���m �ҭ��ǵ;�oN�s������Ʈ��eC�L��L~׭;��O>ի�}�8��lm��r�0A�R ��=�"��<���u��0�需F��1�0� 9�X
 �S����Ú)\Ȝu/YPH�L �8ZK&�A�	!qo�$���f'a��=}>�@�1�qN�r֥_[��1��2F_���P���J�H"	�����8.��_��m�]gs�ö����խ�&oU����UwE%�ʠ���G�M}wR}pa�d��e�,;���~[�A[/U�<��t�*�iW���g߃\ͪl'GU���q���i\�`��'Z���9J�n^u��״nBfkn���&CLJ��p�2J3d���u��L�U��ȰC+a\�2)��4�Zhl��K0ް�ӻK�p���1����3��R�Hѣn����j���]_B��h�	�/d��P��/�_.Ft�ҍ��C�Ov�pk!����ߏ�䩱�??�<�������,U4���wv0����.��b�M�����A�I�+�HNq��܏�oStn
b$E�9b9N�&L BS�5��,���H��͉a�K%毶%_\~�l��6�e�a8�����1E�0�2#�f���]���9(	��e#�R��2��BYir��"�w�r�5ԤA�(bܖ�[HK2nMn�$d�Rt��ʫ����O���ȼJ�p���q"L0F���KL�������J�;�K~=� 6�b]�P�x��?PK
   �I�XX:B�]  �h                  cirkitFile.jsonPK
   �I�X�H<�'  �'  /             �  images/289c84f5-bee9-42dc-8a56-be82ea7098c8.pngPK
   �I�X�ޗԊ  �  /             d?  images/290f8d32-1f39-4e19-80b6-a4526aa84625.pngPK
   oI�X�<0*r�  �
 /             ;P  images/46ec3c75-1d43-4a14-938d-e2b5ecdc5822.jpgPK
   �I�X}�� � /             � images/5874d651-dcf0-4a98-b8b4-9fcbfdf83d7f.pngPK
   x��X?�-�,�  )�  /             0� images/6217b039-096c-42ca-9a04-ba011aa6a0cd.pngPK
   oI�Xډ�'��   �  /             �� images/9b01e4e0-397a-41ff-a8da-0d69e8cd9d76.jpgPK
   x��X`"�v�  ��  /             �p images/adcf2c83-f38d-4d07-a246-237caa0514e4.pngPK
   �I�X�{9� �, /             `_	 images/c24ad21a-d149-4590-811d-5086112a7898.pngPK
   �I�X
V+c  �               �A jsons/user_defined.jsonPK    
 
 j  #H   